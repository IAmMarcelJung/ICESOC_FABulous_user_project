module eFPGA_top
    #(
        parameter include_eFPGA=1,
        parameter NumberOfRows=14,
        parameter NumberOfCols=15,
        parameter FrameBitsPerRow=32,
        parameter MaxFramesPerCol=20,
        parameter desync_flag=20,
        parameter FrameSelectWidth=5,
        parameter RowSelectWidth=5
    )
    (
        //External IO port
        output [19:0] A_config_C,
        output [19:0] B_config_C,
        output [19:0] Config_accessC,
        output [9:0] I_top,
        input [9:0] O_top,
        input [36-1:0] W_OPA,
        input [36-1:0] W_OPB,
        output [36-1:0] W_RES0,
        output [36-1:0] W_RES1,
        output [36-1:0] W_RES2,

        input [36-1:0] E_OPA,
        input [36-1:0] E_OPB,
        output [36-1:0] E_RES0,
        output [36-1:0] E_RES1,
        output [36-1:0] E_RES2,
        output [9:0] T_top,
        //Config related ports
        input CLK,
        input resetn,
        input SelfWriteStrobe,
        input [31:0] SelfWriteData,
        input Rx,
        output ComActive,
        output ReceiveLED,
        input s_clk,
        input s_data
);
 //BlockRAM ports

// /*
// wire[224-1:0] RAM2FAB_D_I;
// wire[224-1:0] FAB2RAM_D_O;
// wire[112-1:0] FAB2RAM_A_O;
// wire[56-1:0] FAB2RAM_C_O;
// */

wire [80-1:0] RAM2FAB_D;
wire [80-1:0] FAB2RAM_D;
wire [40-1:0] FAB2RAM_A;
wire [20-1:0] FAB2RAM_C;

 //Signal declarations
wire[(NumberOfRows*FrameBitsPerRow)-1:0] FrameRegister;
wire[(MaxFramesPerCol*NumberOfCols)-1:0] FrameSelect;
wire[(FrameBitsPerRow*(NumberOfRows+2))-1:0] FrameData;
wire[FrameBitsPerRow-1:0] FrameAddressRegister;
wire LongFrameStrobe;
wire[31:0] LocalWriteData;
wire LocalWriteStrobe;
wire[RowSelectWidth-1:0] RowSelect;
wire resten;
`ifndef EMULATION

eFPGA_Config
    #(
    .RowSelectWidth(RowSelectWidth),
    .NumberOfRows(NumberOfRows),
    .desync_flag(desync_flag),
    .FrameBitsPerRow(FrameBitsPerRow)
    )
    eFPGA_Config_inst
    (
    .CLK(CLK),
    .resetn(resetn),
    .Rx(Rx),
    .ComActive(ComActive),
    .ReceiveLED(ReceiveLED),
    .s_clk(s_clk),
    .s_data(s_data),
    .SelfWriteData(SelfWriteData),
    .SelfWriteStrobe(SelfWriteStrobe),
    .ConfigWriteData(LocalWriteData),
    .ConfigWriteStrobe(LocalWriteStrobe),
    .FrameAddressRegister(FrameAddressRegister),
    .LongFrameStrobe(LongFrameStrobe),
    .RowSelect(RowSelect)
);


Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(1)
    )
    inst_Frame_Data_Reg_0
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[0*FrameBitsPerRow+FrameBitsPerRow-1:0*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(2)
    )
    inst_Frame_Data_Reg_1
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[1*FrameBitsPerRow+FrameBitsPerRow-1:1*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(3)
    )
    inst_Frame_Data_Reg_2
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[2*FrameBitsPerRow+FrameBitsPerRow-1:2*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(4)
    )
    inst_Frame_Data_Reg_3
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[3*FrameBitsPerRow+FrameBitsPerRow-1:3*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(5)
    )
    inst_Frame_Data_Reg_4
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[4*FrameBitsPerRow+FrameBitsPerRow-1:4*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(6)
    )
    inst_Frame_Data_Reg_5
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[5*FrameBitsPerRow+FrameBitsPerRow-1:5*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(7)
    )
    inst_Frame_Data_Reg_6
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[6*FrameBitsPerRow+FrameBitsPerRow-1:6*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(8)
    )
    inst_Frame_Data_Reg_7
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[7*FrameBitsPerRow+FrameBitsPerRow-1:7*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(9)
    )
    inst_Frame_Data_Reg_8
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[8*FrameBitsPerRow+FrameBitsPerRow-1:8*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(10)
    )
    inst_Frame_Data_Reg_9
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[9*FrameBitsPerRow+FrameBitsPerRow-1:9*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(11)
    )
    inst_Frame_Data_Reg_10
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[10*FrameBitsPerRow+FrameBitsPerRow-1:10*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(12)
    )
    inst_Frame_Data_Reg_11
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[11*FrameBitsPerRow+FrameBitsPerRow-1:11*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(13)
    )
    inst_Frame_Data_Reg_12
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[12*FrameBitsPerRow+FrameBitsPerRow-1:12*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(14)
    )
    inst_Frame_Data_Reg_13
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[13*FrameBitsPerRow+FrameBitsPerRow-1:13*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);


Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(0)
    )
    inst_Frame_Select_0
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[0*MaxFramesPerCol+MaxFramesPerCol-1:0*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(1)
    )
    inst_Frame_Select_1
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[1*MaxFramesPerCol+MaxFramesPerCol-1:1*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(2)
    )
    inst_Frame_Select_2
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[2*MaxFramesPerCol+MaxFramesPerCol-1:2*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(3)
    )
    inst_Frame_Select_3
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[3*MaxFramesPerCol+MaxFramesPerCol-1:3*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(4)
    )
    inst_Frame_Select_4
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[4*MaxFramesPerCol+MaxFramesPerCol-1:4*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(5)
    )
    inst_Frame_Select_5
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[5*MaxFramesPerCol+MaxFramesPerCol-1:5*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(6)
    )
    inst_Frame_Select_6
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[6*MaxFramesPerCol+MaxFramesPerCol-1:6*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(7)
    )
    inst_Frame_Select_7
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[7*MaxFramesPerCol+MaxFramesPerCol-1:7*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(8)
    )
    inst_Frame_Select_8
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[8*MaxFramesPerCol+MaxFramesPerCol-1:8*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(9)
    )
    inst_Frame_Select_9
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[9*MaxFramesPerCol+MaxFramesPerCol-1:9*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(10)
    )
    inst_Frame_Select_10
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[10*MaxFramesPerCol+MaxFramesPerCol-1:10*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(11)
    )
    inst_Frame_Select_11
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[11*MaxFramesPerCol+MaxFramesPerCol-1:11*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(12)
    )
    inst_Frame_Select_12
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[12*MaxFramesPerCol+MaxFramesPerCol-1:12*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(13)
    )
    inst_Frame_Select_13
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[13*MaxFramesPerCol+MaxFramesPerCol-1:13*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(14)
    )
    inst_Frame_Select_14
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[14*MaxFramesPerCol+MaxFramesPerCol-1:14*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);


`endif
 eFPGA Inst_eFPGA(
        .Tile_X0Y10_A_I_top(I_top[9]),
        .Tile_X0Y10_B_I_top(I_top[8]),
        .Tile_X0Y11_A_I_top(I_top[7]),
        .Tile_X0Y11_B_I_top(I_top[6]),
        .Tile_X0Y12_A_I_top(I_top[5]),
        .Tile_X0Y12_B_I_top(I_top[4]),
        .Tile_X0Y13_A_I_top(I_top[3]),
        .Tile_X0Y13_B_I_top(I_top[2]),
        .Tile_X0Y14_A_I_top(I_top[1]),
        .Tile_X0Y14_B_I_top(I_top[0]),

        .Tile_X0Y10_A_T_top(T_top[9]),
        .Tile_X0Y10_B_T_top(T_top[8]),
        .Tile_X0Y11_A_T_top(T_top[7]),
        .Tile_X0Y11_B_T_top(T_top[6]),
        .Tile_X0Y12_A_T_top(T_top[5]),
        .Tile_X0Y12_B_T_top(T_top[4]),
        .Tile_X0Y13_A_T_top(T_top[3]),
        .Tile_X0Y13_B_T_top(T_top[2]),
        .Tile_X0Y14_A_T_top(T_top[1]),
        .Tile_X0Y14_B_T_top(T_top[0]),

        .Tile_X0Y10_A_O_top(O_top[9]),
        .Tile_X0Y10_B_O_top(O_top[8]),
        .Tile_X0Y11_A_O_top(O_top[7]),
        .Tile_X0Y11_B_O_top(O_top[6]),
        .Tile_X0Y12_A_O_top(O_top[5]),
        .Tile_X0Y12_B_O_top(O_top[4]),
        .Tile_X0Y13_A_O_top(O_top[3]),
        .Tile_X0Y13_B_O_top(O_top[2]),
        .Tile_X0Y14_A_O_top(O_top[1]),
        .Tile_X0Y14_B_O_top(O_top[0]),

        .Tile_X0Y10_A_config_C_bit0(A_config_C[19]),
        .Tile_X0Y10_A_config_C_bit1(A_config_C[18]),
        .Tile_X0Y10_A_config_C_bit2(A_config_C[17]),
        .Tile_X0Y10_A_config_C_bit3(A_config_C[16]),
        .Tile_X0Y11_A_config_C_bit0(A_config_C[15]),
        .Tile_X0Y11_A_config_C_bit1(A_config_C[14]),
        .Tile_X0Y11_A_config_C_bit2(A_config_C[13]),
        .Tile_X0Y11_A_config_C_bit3(A_config_C[12]),
        .Tile_X0Y12_A_config_C_bit0(A_config_C[11]),
        .Tile_X0Y12_A_config_C_bit1(A_config_C[10]),
        .Tile_X0Y12_A_config_C_bit2(A_config_C[9]),
        .Tile_X0Y12_A_config_C_bit3(A_config_C[8]),
        .Tile_X0Y13_A_config_C_bit0(A_config_C[7]),
        .Tile_X0Y13_A_config_C_bit1(A_config_C[6]),
        .Tile_X0Y13_A_config_C_bit2(A_config_C[5]),
        .Tile_X0Y13_A_config_C_bit3(A_config_C[4]),
        .Tile_X0Y14_A_config_C_bit0(A_config_C[3]),
        .Tile_X0Y14_A_config_C_bit1(A_config_C[2]),
        .Tile_X0Y14_A_config_C_bit2(A_config_C[1]),
        .Tile_X0Y14_A_config_C_bit3(A_config_C[0]),

        .Tile_X0Y10_B_config_C_bit0(B_config_C[19]),
        .Tile_X0Y10_B_config_C_bit1(B_config_C[18]),
        .Tile_X0Y10_B_config_C_bit2(B_config_C[17]),
        .Tile_X0Y10_B_config_C_bit3(B_config_C[16]),
        .Tile_X0Y11_B_config_C_bit0(B_config_C[15]),
        .Tile_X0Y11_B_config_C_bit1(B_config_C[14]),
        .Tile_X0Y11_B_config_C_bit2(B_config_C[13]),
        .Tile_X0Y11_B_config_C_bit3(B_config_C[12]),
        .Tile_X0Y12_B_config_C_bit0(B_config_C[11]),
        .Tile_X0Y12_B_config_C_bit1(B_config_C[10]),
        .Tile_X0Y12_B_config_C_bit2(B_config_C[9]),
        .Tile_X0Y12_B_config_C_bit3(B_config_C[8]),
        .Tile_X0Y13_B_config_C_bit0(B_config_C[7]),
        .Tile_X0Y13_B_config_C_bit1(B_config_C[6]),
        .Tile_X0Y13_B_config_C_bit2(B_config_C[5]),
        .Tile_X0Y13_B_config_C_bit3(B_config_C[4]),
        .Tile_X0Y14_B_config_C_bit0(B_config_C[3]),
        .Tile_X0Y14_B_config_C_bit1(B_config_C[2]),
        .Tile_X0Y14_B_config_C_bit2(B_config_C[1]),
        .Tile_X0Y14_B_config_C_bit3(B_config_C[0]),

        .Tile_X3Y1_OPA_I0(W_OPA[35]),
        .Tile_X3Y1_OPA_I1(W_OPA[34]),
        .Tile_X3Y1_OPA_I2(W_OPA[33]),
        .Tile_X3Y1_OPA_I3(W_OPA[32]),
        .Tile_X3Y2_OPA_I0(W_OPA[31]),
        .Tile_X3Y2_OPA_I1(W_OPA[30]),
        .Tile_X3Y2_OPA_I2(W_OPA[29]),
        .Tile_X3Y2_OPA_I3(W_OPA[28]),
        .Tile_X3Y3_OPA_I0(W_OPA[27]),
        .Tile_X3Y3_OPA_I1(W_OPA[26]),
        .Tile_X3Y3_OPA_I2(W_OPA[25]),
        .Tile_X3Y3_OPA_I3(W_OPA[24]),
        .Tile_X3Y4_OPA_I0(W_OPA[23]),
        .Tile_X3Y4_OPA_I1(W_OPA[22]),
        .Tile_X3Y4_OPA_I2(W_OPA[21]),
        .Tile_X3Y4_OPA_I3(W_OPA[20]),
        .Tile_X3Y5_OPA_I0(W_OPA[19]),
        .Tile_X3Y5_OPA_I1(W_OPA[18]),
        .Tile_X3Y5_OPA_I2(W_OPA[17]),
        .Tile_X3Y5_OPA_I3(W_OPA[16]),
        .Tile_X3Y6_OPA_I0(W_OPA[15]),
        .Tile_X3Y6_OPA_I1(W_OPA[14]),
        .Tile_X3Y6_OPA_I2(W_OPA[13]),
        .Tile_X3Y6_OPA_I3(W_OPA[12]),
        .Tile_X3Y7_OPA_I0(W_OPA[11]),
        .Tile_X3Y7_OPA_I1(W_OPA[10]),
        .Tile_X3Y7_OPA_I2(W_OPA[9]),
        .Tile_X3Y7_OPA_I3(W_OPA[8]),
        .Tile_X3Y8_OPA_I0(W_OPA[7]),
        .Tile_X3Y8_OPA_I1(W_OPA[6]),
        .Tile_X3Y8_OPA_I2(W_OPA[5]),
        .Tile_X3Y8_OPA_I3(W_OPA[4]),
        .Tile_X3Y9_OPA_I0(W_OPA[3]),
        .Tile_X3Y9_OPA_I1(W_OPA[2]),
        .Tile_X3Y9_OPA_I2(W_OPA[1]),
        .Tile_X3Y9_OPA_I3(W_OPA[0]),

        .Tile_X3Y1_OPB_I0(W_OPB[35]),
        .Tile_X3Y1_OPB_I1(W_OPB[34]),
        .Tile_X3Y1_OPB_I2(W_OPB[33]),
        .Tile_X3Y1_OPB_I3(W_OPB[32]),
        .Tile_X3Y2_OPB_I0(W_OPB[31]),
        .Tile_X3Y2_OPB_I1(W_OPB[30]),
        .Tile_X3Y2_OPB_I2(W_OPB[29]),
        .Tile_X3Y2_OPB_I3(W_OPB[28]),
        .Tile_X3Y3_OPB_I0(W_OPB[27]),
        .Tile_X3Y3_OPB_I1(W_OPB[26]),
        .Tile_X3Y3_OPB_I2(W_OPB[25]),
        .Tile_X3Y3_OPB_I3(W_OPB[24]),
        .Tile_X3Y4_OPB_I0(W_OPB[23]),
        .Tile_X3Y4_OPB_I1(W_OPB[22]),
        .Tile_X3Y4_OPB_I2(W_OPB[21]),
        .Tile_X3Y4_OPB_I3(W_OPB[20]),
        .Tile_X3Y5_OPB_I0(W_OPB[19]),
        .Tile_X3Y5_OPB_I1(W_OPB[18]),
        .Tile_X3Y5_OPB_I2(W_OPB[17]),
        .Tile_X3Y5_OPB_I3(W_OPB[16]),
        .Tile_X3Y6_OPB_I0(W_OPB[15]),
        .Tile_X3Y6_OPB_I1(W_OPB[14]),
        .Tile_X3Y6_OPB_I2(W_OPB[13]),
        .Tile_X3Y6_OPB_I3(W_OPB[12]),
        .Tile_X3Y7_OPB_I0(W_OPB[11]),
        .Tile_X3Y7_OPB_I1(W_OPB[10]),
        .Tile_X3Y7_OPB_I2(W_OPB[9]),
        .Tile_X3Y7_OPB_I3(W_OPB[8]),
        .Tile_X3Y8_OPB_I0(W_OPB[7]),
        .Tile_X3Y8_OPB_I1(W_OPB[6]),
        .Tile_X3Y8_OPB_I2(W_OPB[5]),
        .Tile_X3Y8_OPB_I3(W_OPB[4]),
        .Tile_X3Y9_OPB_I0(W_OPB[3]),
        .Tile_X3Y9_OPB_I1(W_OPB[2]),
        .Tile_X3Y9_OPB_I2(W_OPB[1]),
        .Tile_X3Y9_OPB_I3(W_OPB[0]),

        .Tile_X3Y1_RES0_O0(W_RES0[35]),
        .Tile_X3Y1_RES0_O1(W_RES0[34]),
        .Tile_X3Y1_RES0_O2(W_RES0[33]),
        .Tile_X3Y1_RES0_O3(W_RES0[32]),
        .Tile_X3Y2_RES0_O0(W_RES0[31]),
        .Tile_X3Y2_RES0_O1(W_RES0[30]),
        .Tile_X3Y2_RES0_O2(W_RES0[29]),
        .Tile_X3Y2_RES0_O3(W_RES0[28]),
        .Tile_X3Y3_RES0_O0(W_RES0[27]),
        .Tile_X3Y3_RES0_O1(W_RES0[26]),
        .Tile_X3Y3_RES0_O2(W_RES0[25]),
        .Tile_X3Y3_RES0_O3(W_RES0[24]),
        .Tile_X3Y4_RES0_O0(W_RES0[23]),
        .Tile_X3Y4_RES0_O1(W_RES0[22]),
        .Tile_X3Y4_RES0_O2(W_RES0[21]),
        .Tile_X3Y4_RES0_O3(W_RES0[20]),
        .Tile_X3Y5_RES0_O0(W_RES0[19]),
        .Tile_X3Y5_RES0_O1(W_RES0[18]),
        .Tile_X3Y5_RES0_O2(W_RES0[17]),
        .Tile_X3Y5_RES0_O3(W_RES0[16]),
        .Tile_X3Y6_RES0_O0(W_RES0[15]),
        .Tile_X3Y6_RES0_O1(W_RES0[14]),
        .Tile_X3Y6_RES0_O2(W_RES0[13]),
        .Tile_X3Y6_RES0_O3(W_RES0[12]),
        .Tile_X3Y7_RES0_O0(W_RES0[11]),
        .Tile_X3Y7_RES0_O1(W_RES0[10]),
        .Tile_X3Y7_RES0_O2(W_RES0[9]),
        .Tile_X3Y7_RES0_O3(W_RES0[8]),
        .Tile_X3Y8_RES0_O0(W_RES0[7]),
        .Tile_X3Y8_RES0_O1(W_RES0[6]),
        .Tile_X3Y8_RES0_O2(W_RES0[5]),
        .Tile_X3Y8_RES0_O3(W_RES0[4]),
        .Tile_X3Y9_RES0_O0(W_RES0[3]),
        .Tile_X3Y9_RES0_O1(W_RES0[2]),
        .Tile_X3Y9_RES0_O2(W_RES0[1]),
        .Tile_X3Y9_RES0_O3(W_RES0[0]),
	
        .Tile_X3Y1_RES1_O0(W_RES1[35]),
        .Tile_X3Y1_RES1_O1(W_RES1[34]),
        .Tile_X3Y1_RES1_O2(W_RES1[33]),
        .Tile_X3Y1_RES1_O3(W_RES1[32]),
        .Tile_X3Y2_RES1_O0(W_RES1[31]),
        .Tile_X3Y2_RES1_O1(W_RES1[30]),
        .Tile_X3Y2_RES1_O2(W_RES1[29]),
        .Tile_X3Y2_RES1_O3(W_RES1[28]),
        .Tile_X3Y3_RES1_O0(W_RES1[27]),
        .Tile_X3Y3_RES1_O1(W_RES1[26]),
        .Tile_X3Y3_RES1_O2(W_RES1[25]),
        .Tile_X3Y3_RES1_O3(W_RES1[24]),
        .Tile_X3Y4_RES1_O0(W_RES1[23]),
        .Tile_X3Y4_RES1_O1(W_RES1[22]),
        .Tile_X3Y4_RES1_O2(W_RES1[21]),
        .Tile_X3Y4_RES1_O3(W_RES1[20]),
        .Tile_X3Y5_RES1_O0(W_RES1[19]),
        .Tile_X3Y5_RES1_O1(W_RES1[18]),
        .Tile_X3Y5_RES1_O2(W_RES1[17]),
        .Tile_X3Y5_RES1_O3(W_RES1[16]),
        .Tile_X3Y6_RES1_O0(W_RES1[15]),
        .Tile_X3Y6_RES1_O1(W_RES1[14]),
        .Tile_X3Y6_RES1_O2(W_RES1[13]),
        .Tile_X3Y6_RES1_O3(W_RES1[12]),
        .Tile_X3Y7_RES1_O0(W_RES1[11]),
        .Tile_X3Y7_RES1_O1(W_RES1[10]),
        .Tile_X3Y7_RES1_O2(W_RES1[9]),
        .Tile_X3Y7_RES1_O3(W_RES1[8]),
        .Tile_X3Y8_RES1_O0(W_RES1[7]),
        .Tile_X3Y8_RES1_O1(W_RES1[6]),
        .Tile_X3Y8_RES1_O2(W_RES1[5]),
        .Tile_X3Y8_RES1_O3(W_RES1[4]),
        .Tile_X3Y9_RES1_O0(W_RES1[3]),
        .Tile_X3Y9_RES1_O1(W_RES1[2]),
        .Tile_X3Y9_RES1_O2(W_RES1[1]),
        .Tile_X3Y9_RES1_O3(W_RES1[0]),
	
        .Tile_X3Y1_RES2_O0(W_RES2[35]),
        .Tile_X3Y1_RES2_O1(W_RES2[34]),
        .Tile_X3Y1_RES2_O2(W_RES2[33]),
        .Tile_X3Y1_RES2_O3(W_RES2[32]),
        .Tile_X3Y2_RES2_O0(W_RES2[31]),
        .Tile_X3Y2_RES2_O1(W_RES2[30]),
        .Tile_X3Y2_RES2_O2(W_RES2[29]),
        .Tile_X3Y2_RES2_O3(W_RES2[28]),
        .Tile_X3Y3_RES2_O0(W_RES2[27]),
        .Tile_X3Y3_RES2_O1(W_RES2[26]),
        .Tile_X3Y3_RES2_O2(W_RES2[25]),
        .Tile_X3Y3_RES2_O3(W_RES2[24]),
        .Tile_X3Y4_RES2_O0(W_RES2[23]),
        .Tile_X3Y4_RES2_O1(W_RES2[22]),
        .Tile_X3Y4_RES2_O2(W_RES2[21]),
        .Tile_X3Y4_RES2_O3(W_RES2[20]),
        .Tile_X3Y5_RES2_O0(W_RES2[19]),
        .Tile_X3Y5_RES2_O1(W_RES2[18]),
        .Tile_X3Y5_RES2_O2(W_RES2[17]),
        .Tile_X3Y5_RES2_O3(W_RES2[16]),
        .Tile_X3Y6_RES2_O0(W_RES2[15]),
        .Tile_X3Y6_RES2_O1(W_RES2[14]),
        .Tile_X3Y6_RES2_O2(W_RES2[13]),
        .Tile_X3Y6_RES2_O3(W_RES2[12]),
        .Tile_X3Y7_RES2_O0(W_RES2[11]),
        .Tile_X3Y7_RES2_O1(W_RES2[10]),
        .Tile_X3Y7_RES2_O2(W_RES2[9]),
        .Tile_X3Y7_RES2_O3(W_RES2[8]),
        .Tile_X3Y8_RES2_O0(W_RES2[7]),
        .Tile_X3Y8_RES2_O1(W_RES2[6]),
        .Tile_X3Y8_RES2_O2(W_RES2[5]),
        .Tile_X3Y8_RES2_O3(W_RES2[4]),
        .Tile_X3Y9_RES2_O0(W_RES2[3]),
        .Tile_X3Y9_RES2_O1(W_RES2[2]),
        .Tile_X3Y9_RES2_O2(W_RES2[1]),
        .Tile_X3Y9_RES2_O3(W_RES2[0]),

        .Tile_X11Y1_OPA_I0(E_OPA[35]),
        .Tile_X11Y1_OPA_I1(E_OPA[34]),
        .Tile_X11Y1_OPA_I2(E_OPA[33]),
        .Tile_X11Y1_OPA_I3(E_OPA[32]),
        .Tile_X11Y2_OPA_I0(E_OPA[31]),
        .Tile_X11Y2_OPA_I1(E_OPA[30]),
        .Tile_X11Y2_OPA_I2(E_OPA[29]),
        .Tile_X11Y2_OPA_I3(E_OPA[28]),
        .Tile_X11Y3_OPA_I0(E_OPA[27]),
        .Tile_X11Y3_OPA_I1(E_OPA[26]),
        .Tile_X11Y3_OPA_I2(E_OPA[25]),
        .Tile_X11Y3_OPA_I3(E_OPA[24]),
        .Tile_X11Y4_OPA_I0(E_OPA[23]),
        .Tile_X11Y4_OPA_I1(E_OPA[22]),
        .Tile_X11Y4_OPA_I2(E_OPA[21]),
        .Tile_X11Y4_OPA_I3(E_OPA[20]),
        .Tile_X11Y5_OPA_I0(E_OPA[19]),
        .Tile_X11Y5_OPA_I1(E_OPA[18]),
        .Tile_X11Y5_OPA_I2(E_OPA[17]),
        .Tile_X11Y5_OPA_I3(E_OPA[16]),
        .Tile_X11Y6_OPA_I0(E_OPA[15]),
        .Tile_X11Y6_OPA_I1(E_OPA[14]),
        .Tile_X11Y6_OPA_I2(E_OPA[13]),
        .Tile_X11Y6_OPA_I3(E_OPA[12]),
        .Tile_X11Y7_OPA_I0(E_OPA[11]),
        .Tile_X11Y7_OPA_I1(E_OPA[10]),
        .Tile_X11Y7_OPA_I2(E_OPA[9]),
        .Tile_X11Y7_OPA_I3(E_OPA[8]),
        .Tile_X11Y8_OPA_I0(E_OPA[7]),
        .Tile_X11Y8_OPA_I1(E_OPA[6]),
        .Tile_X11Y8_OPA_I2(E_OPA[5]),
        .Tile_X11Y8_OPA_I3(E_OPA[4]),
        .Tile_X11Y9_OPA_I0(E_OPA[3]),
        .Tile_X11Y9_OPA_I1(E_OPA[2]),
        .Tile_X11Y9_OPA_I2(E_OPA[1]),
        .Tile_X11Y9_OPA_I3(E_OPA[0]),
	
        .Tile_X11Y1_OPB_I0(E_OPB[35]),
        .Tile_X11Y1_OPB_I1(E_OPB[34]),
        .Tile_X11Y1_OPB_I2(E_OPB[33]),
        .Tile_X11Y1_OPB_I3(E_OPB[32]),
        .Tile_X11Y2_OPB_I0(E_OPB[31]),
        .Tile_X11Y2_OPB_I1(E_OPB[30]),
        .Tile_X11Y2_OPB_I2(E_OPB[29]),
        .Tile_X11Y2_OPB_I3(E_OPB[28]),
        .Tile_X11Y3_OPB_I0(E_OPB[27]),
        .Tile_X11Y3_OPB_I1(E_OPB[26]),
        .Tile_X11Y3_OPB_I2(E_OPB[25]),
        .Tile_X11Y3_OPB_I3(E_OPB[24]),
        .Tile_X11Y4_OPB_I0(E_OPB[23]),
        .Tile_X11Y4_OPB_I1(E_OPB[22]),
        .Tile_X11Y4_OPB_I2(E_OPB[21]),
        .Tile_X11Y4_OPB_I3(E_OPB[20]),
        .Tile_X11Y5_OPB_I0(E_OPB[19]),
        .Tile_X11Y5_OPB_I1(E_OPB[18]),
        .Tile_X11Y5_OPB_I2(E_OPB[17]),
        .Tile_X11Y5_OPB_I3(E_OPB[16]),
        .Tile_X11Y6_OPB_I0(E_OPB[15]),
        .Tile_X11Y6_OPB_I1(E_OPB[14]),
        .Tile_X11Y6_OPB_I2(E_OPB[13]),
        .Tile_X11Y6_OPB_I3(E_OPB[12]),
        .Tile_X11Y7_OPB_I0(E_OPB[11]),
        .Tile_X11Y7_OPB_I1(E_OPB[10]),
        .Tile_X11Y7_OPB_I2(E_OPB[9]),
        .Tile_X11Y7_OPB_I3(E_OPB[8]),
        .Tile_X11Y8_OPB_I0(E_OPB[7]),
        .Tile_X11Y8_OPB_I1(E_OPB[6]),
        .Tile_X11Y8_OPB_I2(E_OPB[5]),
        .Tile_X11Y8_OPB_I3(E_OPB[4]),
        .Tile_X11Y9_OPB_I0(E_OPB[3]),
        .Tile_X11Y9_OPB_I1(E_OPB[2]),
        .Tile_X11Y9_OPB_I2(E_OPB[1]),
        .Tile_X11Y9_OPB_I3(E_OPB[0]),
	
        .Tile_X11Y1_RES0_O0(E_RES0[35]),
        .Tile_X11Y1_RES0_O1(E_RES0[34]),
        .Tile_X11Y1_RES0_O2(E_RES0[33]),
        .Tile_X11Y1_RES0_O3(E_RES0[32]),
        .Tile_X11Y2_RES0_O0(E_RES0[31]),
        .Tile_X11Y2_RES0_O1(E_RES0[30]),
        .Tile_X11Y2_RES0_O2(E_RES0[29]),
        .Tile_X11Y2_RES0_O3(E_RES0[28]),
        .Tile_X11Y3_RES0_O0(E_RES0[27]),
        .Tile_X11Y3_RES0_O1(E_RES0[26]),
        .Tile_X11Y3_RES0_O2(E_RES0[25]),
        .Tile_X11Y3_RES0_O3(E_RES0[24]),
        .Tile_X11Y4_RES0_O0(E_RES0[23]),
        .Tile_X11Y4_RES0_O1(E_RES0[22]),
        .Tile_X11Y4_RES0_O2(E_RES0[21]),
        .Tile_X11Y4_RES0_O3(E_RES0[20]),
        .Tile_X11Y5_RES0_O0(E_RES0[19]),
        .Tile_X11Y5_RES0_O1(E_RES0[18]),
        .Tile_X11Y5_RES0_O2(E_RES0[17]),
        .Tile_X11Y5_RES0_O3(E_RES0[16]),
        .Tile_X11Y6_RES0_O0(E_RES0[15]),
        .Tile_X11Y6_RES0_O1(E_RES0[14]),
        .Tile_X11Y6_RES0_O2(E_RES0[13]),
        .Tile_X11Y6_RES0_O3(E_RES0[12]),
        .Tile_X11Y7_RES0_O0(E_RES0[11]),
        .Tile_X11Y7_RES0_O1(E_RES0[10]),
        .Tile_X11Y7_RES0_O2(E_RES0[9]),
        .Tile_X11Y7_RES0_O3(E_RES0[8]),
        .Tile_X11Y8_RES0_O0(E_RES0[7]),
        .Tile_X11Y8_RES0_O1(E_RES0[6]),
        .Tile_X11Y8_RES0_O2(E_RES0[5]),
        .Tile_X11Y8_RES0_O3(E_RES0[4]),
        .Tile_X11Y9_RES0_O0(E_RES0[3]),
        .Tile_X11Y9_RES0_O1(E_RES0[2]),
        .Tile_X11Y9_RES0_O2(E_RES0[1]),
        .Tile_X11Y9_RES0_O3(E_RES0[0]),
	
        .Tile_X11Y1_RES1_O0(E_RES1[35]),
        .Tile_X11Y1_RES1_O1(E_RES1[34]),
        .Tile_X11Y1_RES1_O2(E_RES1[33]),
        .Tile_X11Y1_RES1_O3(E_RES1[32]),
        .Tile_X11Y2_RES1_O0(E_RES1[31]),
        .Tile_X11Y2_RES1_O1(E_RES1[30]),
        .Tile_X11Y2_RES1_O2(E_RES1[29]),
        .Tile_X11Y2_RES1_O3(E_RES1[28]),
        .Tile_X11Y3_RES1_O0(E_RES1[27]),
        .Tile_X11Y3_RES1_O1(E_RES1[26]),
        .Tile_X11Y3_RES1_O2(E_RES1[25]),
        .Tile_X11Y3_RES1_O3(E_RES1[24]),
        .Tile_X11Y4_RES1_O0(E_RES1[23]),
        .Tile_X11Y4_RES1_O1(E_RES1[22]),
        .Tile_X11Y4_RES1_O2(E_RES1[21]),
        .Tile_X11Y4_RES1_O3(E_RES1[20]),
        .Tile_X11Y5_RES1_O0(E_RES1[19]),
        .Tile_X11Y5_RES1_O1(E_RES1[18]),
        .Tile_X11Y5_RES1_O2(E_RES1[17]),
        .Tile_X11Y5_RES1_O3(E_RES1[16]),
        .Tile_X11Y6_RES1_O0(E_RES1[15]),
        .Tile_X11Y6_RES1_O1(E_RES1[14]),
        .Tile_X11Y6_RES1_O2(E_RES1[13]),
        .Tile_X11Y6_RES1_O3(E_RES1[12]),
        .Tile_X11Y7_RES1_O0(E_RES1[11]),
        .Tile_X11Y7_RES1_O1(E_RES1[10]),
        .Tile_X11Y7_RES1_O2(E_RES1[9]),
        .Tile_X11Y7_RES1_O3(E_RES1[8]),
        .Tile_X11Y8_RES1_O0(E_RES1[7]),
        .Tile_X11Y8_RES1_O1(E_RES1[6]),
        .Tile_X11Y8_RES1_O2(E_RES1[5]),
        .Tile_X11Y8_RES1_O3(E_RES1[4]),
        .Tile_X11Y9_RES1_O0(E_RES1[3]),
        .Tile_X11Y9_RES1_O1(E_RES1[2]),
        .Tile_X11Y9_RES1_O2(E_RES1[1]),
        .Tile_X11Y9_RES1_O3(E_RES1[0]),
	
        .Tile_X11Y1_RES2_O0(E_RES2[35]),
        .Tile_X11Y1_RES2_O1(E_RES2[34]),
        .Tile_X11Y1_RES2_O2(E_RES2[33]),
        .Tile_X11Y1_RES2_O3(E_RES2[32]),
        .Tile_X11Y2_RES2_O0(E_RES2[31]),
        .Tile_X11Y2_RES2_O1(E_RES2[30]),
        .Tile_X11Y2_RES2_O2(E_RES2[29]),
        .Tile_X11Y2_RES2_O3(E_RES2[28]),
        .Tile_X11Y3_RES2_O0(E_RES2[27]),
        .Tile_X11Y3_RES2_O1(E_RES2[26]),
        .Tile_X11Y3_RES2_O2(E_RES2[25]),
        .Tile_X11Y3_RES2_O3(E_RES2[24]),
        .Tile_X11Y4_RES2_O0(E_RES2[23]),
        .Tile_X11Y4_RES2_O1(E_RES2[22]),
        .Tile_X11Y4_RES2_O2(E_RES2[21]),
        .Tile_X11Y4_RES2_O3(E_RES2[20]),
        .Tile_X11Y5_RES2_O0(E_RES2[19]),
        .Tile_X11Y5_RES2_O1(E_RES2[18]),
        .Tile_X11Y5_RES2_O2(E_RES2[17]),
        .Tile_X11Y5_RES2_O3(E_RES2[16]),
        .Tile_X11Y6_RES2_O0(E_RES2[15]),
        .Tile_X11Y6_RES2_O1(E_RES2[14]),
        .Tile_X11Y6_RES2_O2(E_RES2[13]),
        .Tile_X11Y6_RES2_O3(E_RES2[12]),
        .Tile_X11Y7_RES2_O0(E_RES2[11]),
        .Tile_X11Y7_RES2_O1(E_RES2[10]),
        .Tile_X11Y7_RES2_O2(E_RES2[9]),
        .Tile_X11Y7_RES2_O3(E_RES2[8]),
        .Tile_X11Y8_RES2_O0(E_RES2[7]),
        .Tile_X11Y8_RES2_O1(E_RES2[6]),
        .Tile_X11Y8_RES2_O2(E_RES2[5]),
        .Tile_X11Y8_RES2_O3(E_RES2[4]),
        .Tile_X11Y9_RES2_O0(E_RES2[3]),
        .Tile_X11Y9_RES2_O1(E_RES2[2]),
        .Tile_X11Y9_RES2_O2(E_RES2[1]),
        .Tile_X11Y9_RES2_O3(E_RES2[0]),

        .Tile_X14Y10_RAM2FAB_D0_I0(RAM2FAB_D[79]),
        .Tile_X14Y10_RAM2FAB_D0_I1(RAM2FAB_D[78]),
        .Tile_X14Y10_RAM2FAB_D0_I2(RAM2FAB_D[77]),
        .Tile_X14Y10_RAM2FAB_D0_I3(RAM2FAB_D[76]),
        .Tile_X14Y10_RAM2FAB_D1_I0(RAM2FAB_D[75]),
        .Tile_X14Y10_RAM2FAB_D1_I1(RAM2FAB_D[74]),
        .Tile_X14Y10_RAM2FAB_D1_I2(RAM2FAB_D[73]),
        .Tile_X14Y10_RAM2FAB_D1_I3(RAM2FAB_D[72]),
        .Tile_X14Y10_RAM2FAB_D2_I0(RAM2FAB_D[71]),
        .Tile_X14Y10_RAM2FAB_D2_I1(RAM2FAB_D[70]),
        .Tile_X14Y10_RAM2FAB_D2_I2(RAM2FAB_D[69]),
        .Tile_X14Y10_RAM2FAB_D2_I3(RAM2FAB_D[68]),
        .Tile_X14Y10_RAM2FAB_D3_I0(RAM2FAB_D[67]),
        .Tile_X14Y10_RAM2FAB_D3_I1(RAM2FAB_D[66]),
        .Tile_X14Y10_RAM2FAB_D3_I2(RAM2FAB_D[65]),
        .Tile_X14Y10_RAM2FAB_D3_I3(RAM2FAB_D[64]),
        .Tile_X14Y11_RAM2FAB_D0_I0(RAM2FAB_D[63]),
        .Tile_X14Y11_RAM2FAB_D0_I1(RAM2FAB_D[62]),
        .Tile_X14Y11_RAM2FAB_D0_I2(RAM2FAB_D[61]),
        .Tile_X14Y11_RAM2FAB_D0_I3(RAM2FAB_D[60]),
        .Tile_X14Y11_RAM2FAB_D1_I0(RAM2FAB_D[59]),
        .Tile_X14Y11_RAM2FAB_D1_I1(RAM2FAB_D[58]),
        .Tile_X14Y11_RAM2FAB_D1_I2(RAM2FAB_D[57]),
        .Tile_X14Y11_RAM2FAB_D1_I3(RAM2FAB_D[56]),
        .Tile_X14Y11_RAM2FAB_D2_I0(RAM2FAB_D[55]),
        .Tile_X14Y11_RAM2FAB_D2_I1(RAM2FAB_D[54]),
        .Tile_X14Y11_RAM2FAB_D2_I2(RAM2FAB_D[53]),
        .Tile_X14Y11_RAM2FAB_D2_I3(RAM2FAB_D[52]),
        .Tile_X14Y11_RAM2FAB_D3_I0(RAM2FAB_D[51]),
        .Tile_X14Y11_RAM2FAB_D3_I1(RAM2FAB_D[50]),
        .Tile_X14Y11_RAM2FAB_D3_I2(RAM2FAB_D[49]),
        .Tile_X14Y11_RAM2FAB_D3_I3(RAM2FAB_D[48]),
        .Tile_X14Y12_RAM2FAB_D0_I0(RAM2FAB_D[47]),
        .Tile_X14Y12_RAM2FAB_D0_I1(RAM2FAB_D[46]),
        .Tile_X14Y12_RAM2FAB_D0_I2(RAM2FAB_D[45]),
        .Tile_X14Y12_RAM2FAB_D0_I3(RAM2FAB_D[44]),
        .Tile_X14Y12_RAM2FAB_D1_I0(RAM2FAB_D[43]),
        .Tile_X14Y12_RAM2FAB_D1_I1(RAM2FAB_D[42]),
        .Tile_X14Y12_RAM2FAB_D1_I2(RAM2FAB_D[41]),
        .Tile_X14Y12_RAM2FAB_D1_I3(RAM2FAB_D[40]),
        .Tile_X14Y12_RAM2FAB_D2_I0(RAM2FAB_D[39]),
        .Tile_X14Y12_RAM2FAB_D2_I1(RAM2FAB_D[38]),
        .Tile_X14Y12_RAM2FAB_D2_I2(RAM2FAB_D[37]),
        .Tile_X14Y12_RAM2FAB_D2_I3(RAM2FAB_D[36]),
        .Tile_X14Y12_RAM2FAB_D3_I0(RAM2FAB_D[35]),
        .Tile_X14Y12_RAM2FAB_D3_I1(RAM2FAB_D[34]),
        .Tile_X14Y12_RAM2FAB_D3_I2(RAM2FAB_D[33]),
        .Tile_X14Y12_RAM2FAB_D3_I3(RAM2FAB_D[32]),
        .Tile_X14Y13_RAM2FAB_D0_I0(RAM2FAB_D[31]),
        .Tile_X14Y13_RAM2FAB_D0_I1(RAM2FAB_D[30]),
        .Tile_X14Y13_RAM2FAB_D0_I2(RAM2FAB_D[29]),
        .Tile_X14Y13_RAM2FAB_D0_I3(RAM2FAB_D[28]),
        .Tile_X14Y13_RAM2FAB_D1_I0(RAM2FAB_D[27]),
        .Tile_X14Y13_RAM2FAB_D1_I1(RAM2FAB_D[26]),
        .Tile_X14Y13_RAM2FAB_D1_I2(RAM2FAB_D[25]),
        .Tile_X14Y13_RAM2FAB_D1_I3(RAM2FAB_D[24]),
        .Tile_X14Y13_RAM2FAB_D2_I0(RAM2FAB_D[23]),
        .Tile_X14Y13_RAM2FAB_D2_I1(RAM2FAB_D[22]),
        .Tile_X14Y13_RAM2FAB_D2_I2(RAM2FAB_D[21]),
        .Tile_X14Y13_RAM2FAB_D2_I3(RAM2FAB_D[20]),
        .Tile_X14Y13_RAM2FAB_D3_I0(RAM2FAB_D[19]),
        .Tile_X14Y13_RAM2FAB_D3_I1(RAM2FAB_D[18]),
        .Tile_X14Y13_RAM2FAB_D3_I2(RAM2FAB_D[17]),
        .Tile_X14Y13_RAM2FAB_D3_I3(RAM2FAB_D[16]),
        .Tile_X14Y14_RAM2FAB_D0_I0(RAM2FAB_D[15]),
        .Tile_X14Y14_RAM2FAB_D0_I1(RAM2FAB_D[14]),
        .Tile_X14Y14_RAM2FAB_D0_I2(RAM2FAB_D[13]),
        .Tile_X14Y14_RAM2FAB_D0_I3(RAM2FAB_D[12]),
        .Tile_X14Y14_RAM2FAB_D1_I0(RAM2FAB_D[11]),
        .Tile_X14Y14_RAM2FAB_D1_I1(RAM2FAB_D[10]),
        .Tile_X14Y14_RAM2FAB_D1_I2(RAM2FAB_D[9]),
        .Tile_X14Y14_RAM2FAB_D1_I3(RAM2FAB_D[8]),
        .Tile_X14Y14_RAM2FAB_D2_I0(RAM2FAB_D[7]),
        .Tile_X14Y14_RAM2FAB_D2_I1(RAM2FAB_D[6]),
        .Tile_X14Y14_RAM2FAB_D2_I2(RAM2FAB_D[5]),
        .Tile_X14Y14_RAM2FAB_D2_I3(RAM2FAB_D[4]),
        .Tile_X14Y14_RAM2FAB_D3_I0(RAM2FAB_D[3]),
        .Tile_X14Y14_RAM2FAB_D3_I1(RAM2FAB_D[2]),
        .Tile_X14Y14_RAM2FAB_D3_I2(RAM2FAB_D[1]),
        .Tile_X14Y14_RAM2FAB_D3_I3(RAM2FAB_D[0]),

        .Tile_X14Y10_FAB2RAM_D0_O0(FAB2RAM_D[79]),
        .Tile_X14Y10_FAB2RAM_D0_O1(FAB2RAM_D[78]),
        .Tile_X14Y10_FAB2RAM_D0_O2(FAB2RAM_D[77]),
        .Tile_X14Y10_FAB2RAM_D0_O3(FAB2RAM_D[76]),
        .Tile_X14Y10_FAB2RAM_D1_O0(FAB2RAM_D[75]),
        .Tile_X14Y10_FAB2RAM_D1_O1(FAB2RAM_D[74]),
        .Tile_X14Y10_FAB2RAM_D1_O2(FAB2RAM_D[73]),
        .Tile_X14Y10_FAB2RAM_D1_O3(FAB2RAM_D[72]),
        .Tile_X14Y10_FAB2RAM_D2_O0(FAB2RAM_D[71]),
        .Tile_X14Y10_FAB2RAM_D2_O1(FAB2RAM_D[70]),
        .Tile_X14Y10_FAB2RAM_D2_O2(FAB2RAM_D[69]),
        .Tile_X14Y10_FAB2RAM_D2_O3(FAB2RAM_D[68]),
        .Tile_X14Y10_FAB2RAM_D3_O0(FAB2RAM_D[67]),
        .Tile_X14Y10_FAB2RAM_D3_O1(FAB2RAM_D[66]),
        .Tile_X14Y10_FAB2RAM_D3_O2(FAB2RAM_D[65]),
        .Tile_X14Y10_FAB2RAM_D3_O3(FAB2RAM_D[64]),
        .Tile_X14Y11_FAB2RAM_D0_O0(FAB2RAM_D[63]),
        .Tile_X14Y11_FAB2RAM_D0_O1(FAB2RAM_D[62]),
        .Tile_X14Y11_FAB2RAM_D0_O2(FAB2RAM_D[61]),
        .Tile_X14Y11_FAB2RAM_D0_O3(FAB2RAM_D[60]),
        .Tile_X14Y11_FAB2RAM_D1_O0(FAB2RAM_D[59]),
        .Tile_X14Y11_FAB2RAM_D1_O1(FAB2RAM_D[58]),
        .Tile_X14Y11_FAB2RAM_D1_O2(FAB2RAM_D[57]),
        .Tile_X14Y11_FAB2RAM_D1_O3(FAB2RAM_D[56]),
        .Tile_X14Y11_FAB2RAM_D2_O0(FAB2RAM_D[55]),
        .Tile_X14Y11_FAB2RAM_D2_O1(FAB2RAM_D[54]),
        .Tile_X14Y11_FAB2RAM_D2_O2(FAB2RAM_D[53]),
        .Tile_X14Y11_FAB2RAM_D2_O3(FAB2RAM_D[52]),
        .Tile_X14Y11_FAB2RAM_D3_O0(FAB2RAM_D[51]),
        .Tile_X14Y11_FAB2RAM_D3_O1(FAB2RAM_D[50]),
        .Tile_X14Y11_FAB2RAM_D3_O2(FAB2RAM_D[49]),
        .Tile_X14Y11_FAB2RAM_D3_O3(FAB2RAM_D[48]),
        .Tile_X14Y12_FAB2RAM_D0_O0(FAB2RAM_D[47]),
        .Tile_X14Y12_FAB2RAM_D0_O1(FAB2RAM_D[46]),
        .Tile_X14Y12_FAB2RAM_D0_O2(FAB2RAM_D[45]),
        .Tile_X14Y12_FAB2RAM_D0_O3(FAB2RAM_D[44]),
        .Tile_X14Y12_FAB2RAM_D1_O0(FAB2RAM_D[43]),
        .Tile_X14Y12_FAB2RAM_D1_O1(FAB2RAM_D[42]),
        .Tile_X14Y12_FAB2RAM_D1_O2(FAB2RAM_D[41]),
        .Tile_X14Y12_FAB2RAM_D1_O3(FAB2RAM_D[40]),
        .Tile_X14Y12_FAB2RAM_D2_O0(FAB2RAM_D[39]),
        .Tile_X14Y12_FAB2RAM_D2_O1(FAB2RAM_D[38]),
        .Tile_X14Y12_FAB2RAM_D2_O2(FAB2RAM_D[37]),
        .Tile_X14Y12_FAB2RAM_D2_O3(FAB2RAM_D[36]),
        .Tile_X14Y12_FAB2RAM_D3_O0(FAB2RAM_D[35]),
        .Tile_X14Y12_FAB2RAM_D3_O1(FAB2RAM_D[34]),
        .Tile_X14Y12_FAB2RAM_D3_O2(FAB2RAM_D[33]),
        .Tile_X14Y12_FAB2RAM_D3_O3(FAB2RAM_D[32]),
        .Tile_X14Y13_FAB2RAM_D0_O0(FAB2RAM_D[31]),
        .Tile_X14Y13_FAB2RAM_D0_O1(FAB2RAM_D[30]),
        .Tile_X14Y13_FAB2RAM_D0_O2(FAB2RAM_D[29]),
        .Tile_X14Y13_FAB2RAM_D0_O3(FAB2RAM_D[28]),
        .Tile_X14Y13_FAB2RAM_D1_O0(FAB2RAM_D[27]),
        .Tile_X14Y13_FAB2RAM_D1_O1(FAB2RAM_D[26]),
        .Tile_X14Y13_FAB2RAM_D1_O2(FAB2RAM_D[25]),
        .Tile_X14Y13_FAB2RAM_D1_O3(FAB2RAM_D[24]),
        .Tile_X14Y13_FAB2RAM_D2_O0(FAB2RAM_D[23]),
        .Tile_X14Y13_FAB2RAM_D2_O1(FAB2RAM_D[22]),
        .Tile_X14Y13_FAB2RAM_D2_O2(FAB2RAM_D[21]),
        .Tile_X14Y13_FAB2RAM_D2_O3(FAB2RAM_D[20]),
        .Tile_X14Y13_FAB2RAM_D3_O0(FAB2RAM_D[19]),
        .Tile_X14Y13_FAB2RAM_D3_O1(FAB2RAM_D[18]),
        .Tile_X14Y13_FAB2RAM_D3_O2(FAB2RAM_D[17]),
        .Tile_X14Y13_FAB2RAM_D3_O3(FAB2RAM_D[16]),
        .Tile_X14Y14_FAB2RAM_D0_O0(FAB2RAM_D[15]),
        .Tile_X14Y14_FAB2RAM_D0_O1(FAB2RAM_D[14]),
        .Tile_X14Y14_FAB2RAM_D0_O2(FAB2RAM_D[13]),
        .Tile_X14Y14_FAB2RAM_D0_O3(FAB2RAM_D[12]),
        .Tile_X14Y14_FAB2RAM_D1_O0(FAB2RAM_D[11]),
        .Tile_X14Y14_FAB2RAM_D1_O1(FAB2RAM_D[10]),
        .Tile_X14Y14_FAB2RAM_D1_O2(FAB2RAM_D[9]),
        .Tile_X14Y14_FAB2RAM_D1_O3(FAB2RAM_D[8]),
        .Tile_X14Y14_FAB2RAM_D2_O0(FAB2RAM_D[7]),
        .Tile_X14Y14_FAB2RAM_D2_O1(FAB2RAM_D[6]),
        .Tile_X14Y14_FAB2RAM_D2_O2(FAB2RAM_D[5]),
        .Tile_X14Y14_FAB2RAM_D2_O3(FAB2RAM_D[4]),
        .Tile_X14Y14_FAB2RAM_D3_O0(FAB2RAM_D[3]),
        .Tile_X14Y14_FAB2RAM_D3_O1(FAB2RAM_D[2]),
        .Tile_X14Y14_FAB2RAM_D3_O2(FAB2RAM_D[1]),
        .Tile_X14Y14_FAB2RAM_D3_O3(FAB2RAM_D[0]),

        .Tile_X14Y10_FAB2RAM_A0_O0(FAB2RAM_A[39]),
        .Tile_X14Y10_FAB2RAM_A0_O1(FAB2RAM_A[38]),
        .Tile_X14Y10_FAB2RAM_A0_O2(FAB2RAM_A[37]),
        .Tile_X14Y10_FAB2RAM_A0_O3(FAB2RAM_A[36]),
        .Tile_X14Y10_FAB2RAM_A1_O0(FAB2RAM_A[35]),
        .Tile_X14Y10_FAB2RAM_A1_O1(FAB2RAM_A[34]),
        .Tile_X14Y10_FAB2RAM_A1_O2(FAB2RAM_A[33]),
        .Tile_X14Y10_FAB2RAM_A1_O3(FAB2RAM_A[32]),
        .Tile_X14Y11_FAB2RAM_A0_O0(FAB2RAM_A[31]),
        .Tile_X14Y11_FAB2RAM_A0_O1(FAB2RAM_A[30]),
        .Tile_X14Y11_FAB2RAM_A0_O2(FAB2RAM_A[29]),
        .Tile_X14Y11_FAB2RAM_A0_O3(FAB2RAM_A[28]),
        .Tile_X14Y11_FAB2RAM_A1_O0(FAB2RAM_A[27]),
        .Tile_X14Y11_FAB2RAM_A1_O1(FAB2RAM_A[26]),
        .Tile_X14Y11_FAB2RAM_A1_O2(FAB2RAM_A[25]),
        .Tile_X14Y11_FAB2RAM_A1_O3(FAB2RAM_A[24]),
        .Tile_X14Y12_FAB2RAM_A0_O0(FAB2RAM_A[23]),
        .Tile_X14Y12_FAB2RAM_A0_O1(FAB2RAM_A[22]),
        .Tile_X14Y12_FAB2RAM_A0_O2(FAB2RAM_A[21]),
        .Tile_X14Y12_FAB2RAM_A0_O3(FAB2RAM_A[20]),
        .Tile_X14Y12_FAB2RAM_A1_O0(FAB2RAM_A[19]),
        .Tile_X14Y12_FAB2RAM_A1_O1(FAB2RAM_A[18]),
        .Tile_X14Y12_FAB2RAM_A1_O2(FAB2RAM_A[17]),
        .Tile_X14Y12_FAB2RAM_A1_O3(FAB2RAM_A[16]),
        .Tile_X14Y13_FAB2RAM_A0_O0(FAB2RAM_A[15]),
        .Tile_X14Y13_FAB2RAM_A0_O1(FAB2RAM_A[14]),
        .Tile_X14Y13_FAB2RAM_A0_O2(FAB2RAM_A[13]),
        .Tile_X14Y13_FAB2RAM_A0_O3(FAB2RAM_A[12]),
        .Tile_X14Y13_FAB2RAM_A1_O0(FAB2RAM_A[11]),
        .Tile_X14Y13_FAB2RAM_A1_O1(FAB2RAM_A[10]),
        .Tile_X14Y13_FAB2RAM_A1_O2(FAB2RAM_A[9]),
        .Tile_X14Y13_FAB2RAM_A1_O3(FAB2RAM_A[8]),
        .Tile_X14Y14_FAB2RAM_A0_O0(FAB2RAM_A[7]),
        .Tile_X14Y14_FAB2RAM_A0_O1(FAB2RAM_A[6]),
        .Tile_X14Y14_FAB2RAM_A0_O2(FAB2RAM_A[5]),
        .Tile_X14Y14_FAB2RAM_A0_O3(FAB2RAM_A[4]),
        .Tile_X14Y14_FAB2RAM_A1_O0(FAB2RAM_A[3]),
        .Tile_X14Y14_FAB2RAM_A1_O1(FAB2RAM_A[2]),
        .Tile_X14Y14_FAB2RAM_A1_O2(FAB2RAM_A[1]),
        .Tile_X14Y14_FAB2RAM_A1_O3(FAB2RAM_A[0]),

        .Tile_X14Y10_FAB2RAM_C_O0(FAB2RAM_C[19]),
        .Tile_X14Y10_FAB2RAM_C_O1(FAB2RAM_C[18]),
        .Tile_X14Y10_FAB2RAM_C_O2(FAB2RAM_C[17]),
        .Tile_X14Y10_FAB2RAM_C_O3(FAB2RAM_C[16]),
        .Tile_X14Y11_FAB2RAM_C_O0(FAB2RAM_C[15]),
        .Tile_X14Y11_FAB2RAM_C_O1(FAB2RAM_C[14]),
        .Tile_X14Y11_FAB2RAM_C_O2(FAB2RAM_C[13]),
        .Tile_X14Y11_FAB2RAM_C_O3(FAB2RAM_C[12]),
        .Tile_X14Y12_FAB2RAM_C_O0(FAB2RAM_C[11]),
        .Tile_X14Y12_FAB2RAM_C_O1(FAB2RAM_C[10]),
        .Tile_X14Y12_FAB2RAM_C_O2(FAB2RAM_C[9]),
        .Tile_X14Y12_FAB2RAM_C_O3(FAB2RAM_C[8]),
        .Tile_X14Y13_FAB2RAM_C_O0(FAB2RAM_C[7]),
        .Tile_X14Y13_FAB2RAM_C_O1(FAB2RAM_C[6]),
        .Tile_X14Y13_FAB2RAM_C_O2(FAB2RAM_C[5]),
        .Tile_X14Y13_FAB2RAM_C_O3(FAB2RAM_C[4]),
        .Tile_X14Y14_FAB2RAM_C_O0(FAB2RAM_C[3]),
        .Tile_X14Y14_FAB2RAM_C_O1(FAB2RAM_C[2]),
        .Tile_X14Y14_FAB2RAM_C_O2(FAB2RAM_C[1]),
        .Tile_X14Y14_FAB2RAM_C_O3(FAB2RAM_C[0]),

        .Tile_X14Y10_Config_accessC_bit0(Config_accessC[19]),
        .Tile_X14Y10_Config_accessC_bit1(Config_accessC[18]),
        .Tile_X14Y10_Config_accessC_bit2(Config_accessC[17]),
        .Tile_X14Y10_Config_accessC_bit3(Config_accessC[16]),
        .Tile_X14Y11_Config_accessC_bit0(Config_accessC[15]),
        .Tile_X14Y11_Config_accessC_bit1(Config_accessC[14]),
        .Tile_X14Y11_Config_accessC_bit2(Config_accessC[13]),
        .Tile_X14Y11_Config_accessC_bit3(Config_accessC[12]),
        .Tile_X14Y12_Config_accessC_bit0(Config_accessC[11]),
        .Tile_X14Y12_Config_accessC_bit1(Config_accessC[10]),
        .Tile_X14Y12_Config_accessC_bit2(Config_accessC[9]),
        .Tile_X14Y12_Config_accessC_bit3(Config_accessC[8]),
        .Tile_X14Y13_Config_accessC_bit0(Config_accessC[7]),
        .Tile_X14Y13_Config_accessC_bit1(Config_accessC[6]),
        .Tile_X14Y13_Config_accessC_bit2(Config_accessC[5]),
        .Tile_X14Y13_Config_accessC_bit3(Config_accessC[4]),
        .Tile_X14Y14_Config_accessC_bit0(Config_accessC[3]),
        .Tile_X14Y14_Config_accessC_bit1(Config_accessC[2]),
        .Tile_X14Y14_Config_accessC_bit2(Config_accessC[1]),
        .Tile_X14Y14_Config_accessC_bit3(Config_accessC[0]),

        //declarations
        .UserCLK(CLK),
        .FrameData(FrameData),
        .FrameStrobe(FrameSelect)
    );
/*
eFPGA eFPGA_inst (
    .Tile_X0Y14_A_config_C_bit0(A_config_C[0]),
    .Tile_X0Y14_A_config_C_bit1(A_config_C[1]),
    .Tile_X0Y14_A_config_C_bit2(A_config_C[2]),
    .Tile_X0Y14_A_config_C_bit3(A_config_C[3]),
    .Tile_X0Y13_A_config_C_bit0(A_config_C[4]),
    .Tile_X0Y13_A_config_C_bit1(A_config_C[5]),
    .Tile_X0Y13_A_config_C_bit2(A_config_C[6]),
    .Tile_X0Y13_A_config_C_bit3(A_config_C[7]),
    .Tile_X0Y12_A_config_C_bit0(A_config_C[8]),
    .Tile_X0Y12_A_config_C_bit1(A_config_C[9]),
    .Tile_X0Y12_A_config_C_bit2(A_config_C[10]),
    .Tile_X0Y12_A_config_C_bit3(A_config_C[11]),
    .Tile_X0Y11_A_config_C_bit0(A_config_C[12]),
    .Tile_X0Y11_A_config_C_bit1(A_config_C[13]),
    .Tile_X0Y11_A_config_C_bit2(A_config_C[14]),
    .Tile_X0Y11_A_config_C_bit3(A_config_C[15]),
    .Tile_X0Y10_A_config_C_bit0(A_config_C[16]),
    .Tile_X0Y10_A_config_C_bit1(A_config_C[17]),
    .Tile_X0Y10_A_config_C_bit2(A_config_C[18]),
    .Tile_X0Y10_A_config_C_bit3(A_config_C[19]),
    .Tile_X0Y14_B_config_C_bit0(B_config_C[0]),
    .Tile_X0Y14_B_config_C_bit1(B_config_C[1]),
    .Tile_X0Y14_B_config_C_bit2(B_config_C[2]),
    .Tile_X0Y14_B_config_C_bit3(B_config_C[3]),
    .Tile_X0Y13_B_config_C_bit0(B_config_C[4]),
    .Tile_X0Y13_B_config_C_bit1(B_config_C[5]),
    .Tile_X0Y13_B_config_C_bit2(B_config_C[6]),
    .Tile_X0Y13_B_config_C_bit3(B_config_C[7]),
    .Tile_X0Y12_B_config_C_bit0(B_config_C[8]),
    .Tile_X0Y12_B_config_C_bit1(B_config_C[9]),
    .Tile_X0Y12_B_config_C_bit2(B_config_C[10]),
    .Tile_X0Y12_B_config_C_bit3(B_config_C[11]),
    .Tile_X0Y11_B_config_C_bit0(B_config_C[12]),
    .Tile_X0Y11_B_config_C_bit1(B_config_C[13]),
    .Tile_X0Y11_B_config_C_bit2(B_config_C[14]),
    .Tile_X0Y11_B_config_C_bit3(B_config_C[15]),
    .Tile_X0Y10_B_config_C_bit0(B_config_C[16]),
    .Tile_X0Y10_B_config_C_bit1(B_config_C[17]),
    .Tile_X0Y10_B_config_C_bit2(B_config_C[18]),
    .Tile_X0Y10_B_config_C_bit3(B_config_C[19]),
    .Tile_X14Y14_Config_accessC_bit0(Config_accessC[0]),
    .Tile_X14Y14_Config_accessC_bit1(Config_accessC[1]),
    .Tile_X14Y14_Config_accessC_bit2(Config_accessC[2]),
    .Tile_X14Y14_Config_accessC_bit3(Config_accessC[3]),
    .Tile_X14Y13_Config_accessC_bit0(Config_accessC[4]),
    .Tile_X14Y13_Config_accessC_bit1(Config_accessC[5]),
    .Tile_X14Y13_Config_accessC_bit2(Config_accessC[6]),
    .Tile_X14Y13_Config_accessC_bit3(Config_accessC[7]),
    .Tile_X14Y12_Config_accessC_bit0(Config_accessC[8]),
    .Tile_X14Y12_Config_accessC_bit1(Config_accessC[9]),
    .Tile_X14Y12_Config_accessC_bit2(Config_accessC[10]),
    .Tile_X14Y12_Config_accessC_bit3(Config_accessC[11]),
    .Tile_X14Y11_Config_accessC_bit0(Config_accessC[12]),
    .Tile_X14Y11_Config_accessC_bit1(Config_accessC[13]),
    .Tile_X14Y11_Config_accessC_bit2(Config_accessC[14]),
    .Tile_X14Y11_Config_accessC_bit3(Config_accessC[15]),
    .Tile_X14Y10_Config_accessC_bit0(Config_accessC[16]),
    .Tile_X14Y10_Config_accessC_bit1(Config_accessC[17]),
    .Tile_X14Y10_Config_accessC_bit2(Config_accessC[18]),
    .Tile_X14Y10_Config_accessC_bit3(Config_accessC[19]),
    .Tile_X14Y14_FAB2RAM_A0_O0(FAB2RAM_A_O[0]),
    .Tile_X14Y14_FAB2RAM_A0_O1(FAB2RAM_A_O[1]),
    .Tile_X14Y14_FAB2RAM_A0_O2(FAB2RAM_A_O[2]),
    .Tile_X14Y14_FAB2RAM_A0_O3(FAB2RAM_A_O[3]),
    .Tile_X14Y14_FAB2RAM_A1_O0(FAB2RAM_A_O[4]),
    .Tile_X14Y14_FAB2RAM_A1_O1(FAB2RAM_A_O[5]),
    .Tile_X14Y14_FAB2RAM_A1_O2(FAB2RAM_A_O[6]),
    .Tile_X14Y14_FAB2RAM_A1_O3(FAB2RAM_A_O[7]),
    .Tile_X14Y13_FAB2RAM_A0_O0(FAB2RAM_A_O[8]),
    .Tile_X14Y13_FAB2RAM_A0_O1(FAB2RAM_A_O[9]),
    .Tile_X14Y13_FAB2RAM_A0_O2(FAB2RAM_A_O[10]),
    .Tile_X14Y13_FAB2RAM_A0_O3(FAB2RAM_A_O[11]),
    .Tile_X14Y13_FAB2RAM_A1_O0(FAB2RAM_A_O[12]),
    .Tile_X14Y13_FAB2RAM_A1_O1(FAB2RAM_A_O[13]),
    .Tile_X14Y13_FAB2RAM_A1_O2(FAB2RAM_A_O[14]),
    .Tile_X14Y13_FAB2RAM_A1_O3(FAB2RAM_A_O[15]),
    .Tile_X14Y12_FAB2RAM_A0_O0(FAB2RAM_A_O[16]),
    .Tile_X14Y12_FAB2RAM_A0_O1(FAB2RAM_A_O[17]),
    .Tile_X14Y12_FAB2RAM_A0_O2(FAB2RAM_A_O[18]),
    .Tile_X14Y12_FAB2RAM_A0_O3(FAB2RAM_A_O[19]),
    .Tile_X14Y12_FAB2RAM_A1_O0(FAB2RAM_A_O[20]),
    .Tile_X14Y12_FAB2RAM_A1_O1(FAB2RAM_A_O[21]),
    .Tile_X14Y12_FAB2RAM_A1_O2(FAB2RAM_A_O[22]),
    .Tile_X14Y12_FAB2RAM_A1_O3(FAB2RAM_A_O[23]),
    .Tile_X14Y11_FAB2RAM_A0_O0(FAB2RAM_A_O[24]),
    .Tile_X14Y11_FAB2RAM_A0_O1(FAB2RAM_A_O[25]),
    .Tile_X14Y11_FAB2RAM_A0_O2(FAB2RAM_A_O[26]),
    .Tile_X14Y11_FAB2RAM_A0_O3(FAB2RAM_A_O[27]),
    .Tile_X14Y11_FAB2RAM_A1_O0(FAB2RAM_A_O[28]),
    .Tile_X14Y11_FAB2RAM_A1_O1(FAB2RAM_A_O[29]),
    .Tile_X14Y11_FAB2RAM_A1_O2(FAB2RAM_A_O[30]),
    .Tile_X14Y11_FAB2RAM_A1_O3(FAB2RAM_A_O[31]),
    .Tile_X14Y10_FAB2RAM_A0_O0(FAB2RAM_A_O[32]),
    .Tile_X14Y10_FAB2RAM_A0_O1(FAB2RAM_A_O[33]),
    .Tile_X14Y10_FAB2RAM_A0_O2(FAB2RAM_A_O[34]),
    .Tile_X14Y10_FAB2RAM_A0_O3(FAB2RAM_A_O[35]),
    .Tile_X14Y10_FAB2RAM_A1_O0(FAB2RAM_A_O[36]),
    .Tile_X14Y10_FAB2RAM_A1_O1(FAB2RAM_A_O[37]),
    .Tile_X14Y10_FAB2RAM_A1_O2(FAB2RAM_A_O[38]),
    .Tile_X14Y10_FAB2RAM_A1_O3(FAB2RAM_A_O[39]),
    .Tile_X14Y14_FAB2RAM_C_O0(FAB2RAM_C_O[0]),
    .Tile_X14Y14_FAB2RAM_C_O1(FAB2RAM_C_O[1]),
    .Tile_X14Y14_FAB2RAM_C_O2(FAB2RAM_C_O[2]),
    .Tile_X14Y14_FAB2RAM_C_O3(FAB2RAM_C_O[3]),
    .Tile_X14Y13_FAB2RAM_C_O0(FAB2RAM_C_O[4]),
    .Tile_X14Y13_FAB2RAM_C_O1(FAB2RAM_C_O[5]),
    .Tile_X14Y13_FAB2RAM_C_O2(FAB2RAM_C_O[6]),
    .Tile_X14Y13_FAB2RAM_C_O3(FAB2RAM_C_O[7]),
    .Tile_X14Y12_FAB2RAM_C_O0(FAB2RAM_C_O[8]),
    .Tile_X14Y12_FAB2RAM_C_O1(FAB2RAM_C_O[9]),
    .Tile_X14Y12_FAB2RAM_C_O2(FAB2RAM_C_O[10]),
    .Tile_X14Y12_FAB2RAM_C_O3(FAB2RAM_C_O[11]),
    .Tile_X14Y11_FAB2RAM_C_O0(FAB2RAM_C_O[12]),
    .Tile_X14Y11_FAB2RAM_C_O1(FAB2RAM_C_O[13]),
    .Tile_X14Y11_FAB2RAM_C_O2(FAB2RAM_C_O[14]),
    .Tile_X14Y11_FAB2RAM_C_O3(FAB2RAM_C_O[15]),
    .Tile_X14Y10_FAB2RAM_C_O0(FAB2RAM_C_O[16]),
    .Tile_X14Y10_FAB2RAM_C_O1(FAB2RAM_C_O[17]),
    .Tile_X14Y10_FAB2RAM_C_O2(FAB2RAM_C_O[18]),
    .Tile_X14Y10_FAB2RAM_C_O3(FAB2RAM_C_O[19]),
    .Tile_X14Y14_FAB2RAM_D0_O0(FAB2RAM_D_O[0]),
    .Tile_X14Y14_FAB2RAM_D0_O1(FAB2RAM_D_O[1]),
    .Tile_X14Y14_FAB2RAM_D0_O2(FAB2RAM_D_O[2]),
    .Tile_X14Y14_FAB2RAM_D0_O3(FAB2RAM_D_O[3]),
    .Tile_X14Y14_FAB2RAM_D1_O0(FAB2RAM_D_O[4]),
    .Tile_X14Y14_FAB2RAM_D1_O1(FAB2RAM_D_O[5]),
    .Tile_X14Y14_FAB2RAM_D1_O2(FAB2RAM_D_O[6]),
    .Tile_X14Y14_FAB2RAM_D1_O3(FAB2RAM_D_O[7]),
    .Tile_X14Y14_FAB2RAM_D2_O0(FAB2RAM_D_O[8]),
    .Tile_X14Y14_FAB2RAM_D2_O1(FAB2RAM_D_O[9]),
    .Tile_X14Y14_FAB2RAM_D2_O2(FAB2RAM_D_O[10]),
    .Tile_X14Y14_FAB2RAM_D2_O3(FAB2RAM_D_O[11]),
    .Tile_X14Y14_FAB2RAM_D3_O0(FAB2RAM_D_O[12]),
    .Tile_X14Y14_FAB2RAM_D3_O1(FAB2RAM_D_O[13]),
    .Tile_X14Y14_FAB2RAM_D3_O2(FAB2RAM_D_O[14]),
    .Tile_X14Y14_FAB2RAM_D3_O3(FAB2RAM_D_O[15]),
    .Tile_X14Y13_FAB2RAM_D0_O0(FAB2RAM_D_O[16]),
    .Tile_X14Y13_FAB2RAM_D0_O1(FAB2RAM_D_O[17]),
    .Tile_X14Y13_FAB2RAM_D0_O2(FAB2RAM_D_O[18]),
    .Tile_X14Y13_FAB2RAM_D0_O3(FAB2RAM_D_O[19]),
    .Tile_X14Y13_FAB2RAM_D1_O0(FAB2RAM_D_O[20]),
    .Tile_X14Y13_FAB2RAM_D1_O1(FAB2RAM_D_O[21]),
    .Tile_X14Y13_FAB2RAM_D1_O2(FAB2RAM_D_O[22]),
    .Tile_X14Y13_FAB2RAM_D1_O3(FAB2RAM_D_O[23]),
    .Tile_X14Y13_FAB2RAM_D2_O0(FAB2RAM_D_O[24]),
    .Tile_X14Y13_FAB2RAM_D2_O1(FAB2RAM_D_O[25]),
    .Tile_X14Y13_FAB2RAM_D2_O2(FAB2RAM_D_O[26]),
    .Tile_X14Y13_FAB2RAM_D2_O3(FAB2RAM_D_O[27]),
    .Tile_X14Y13_FAB2RAM_D3_O0(FAB2RAM_D_O[28]),
    .Tile_X14Y13_FAB2RAM_D3_O1(FAB2RAM_D_O[29]),
    .Tile_X14Y13_FAB2RAM_D3_O2(FAB2RAM_D_O[30]),
    .Tile_X14Y13_FAB2RAM_D3_O3(FAB2RAM_D_O[31]),
    .Tile_X14Y12_FAB2RAM_D0_O0(FAB2RAM_D_O[32]),
    .Tile_X14Y12_FAB2RAM_D0_O1(FAB2RAM_D_O[33]),
    .Tile_X14Y12_FAB2RAM_D0_O2(FAB2RAM_D_O[34]),
    .Tile_X14Y12_FAB2RAM_D0_O3(FAB2RAM_D_O[35]),
    .Tile_X14Y12_FAB2RAM_D1_O0(FAB2RAM_D_O[36]),
    .Tile_X14Y12_FAB2RAM_D1_O1(FAB2RAM_D_O[37]),
    .Tile_X14Y12_FAB2RAM_D1_O2(FAB2RAM_D_O[38]),
    .Tile_X14Y12_FAB2RAM_D1_O3(FAB2RAM_D_O[39]),
    .Tile_X14Y12_FAB2RAM_D2_O0(FAB2RAM_D_O[40]),
    .Tile_X14Y12_FAB2RAM_D2_O1(FAB2RAM_D_O[41]),
    .Tile_X14Y12_FAB2RAM_D2_O2(FAB2RAM_D_O[42]),
    .Tile_X14Y12_FAB2RAM_D2_O3(FAB2RAM_D_O[43]),
    .Tile_X14Y12_FAB2RAM_D3_O0(FAB2RAM_D_O[44]),
    .Tile_X14Y12_FAB2RAM_D3_O1(FAB2RAM_D_O[45]),
    .Tile_X14Y12_FAB2RAM_D3_O2(FAB2RAM_D_O[46]),
    .Tile_X14Y12_FAB2RAM_D3_O3(FAB2RAM_D_O[47]),
    .Tile_X14Y11_FAB2RAM_D0_O0(FAB2RAM_D_O[48]),
    .Tile_X14Y11_FAB2RAM_D0_O1(FAB2RAM_D_O[49]),
    .Tile_X14Y11_FAB2RAM_D0_O2(FAB2RAM_D_O[50]),
    .Tile_X14Y11_FAB2RAM_D0_O3(FAB2RAM_D_O[51]),
    .Tile_X14Y11_FAB2RAM_D1_O0(FAB2RAM_D_O[52]),
    .Tile_X14Y11_FAB2RAM_D1_O1(FAB2RAM_D_O[53]),
    .Tile_X14Y11_FAB2RAM_D1_O2(FAB2RAM_D_O[54]),
    .Tile_X14Y11_FAB2RAM_D1_O3(FAB2RAM_D_O[55]),
    .Tile_X14Y11_FAB2RAM_D2_O0(FAB2RAM_D_O[56]),
    .Tile_X14Y11_FAB2RAM_D2_O1(FAB2RAM_D_O[57]),
    .Tile_X14Y11_FAB2RAM_D2_O2(FAB2RAM_D_O[58]),
    .Tile_X14Y11_FAB2RAM_D2_O3(FAB2RAM_D_O[59]),
    .Tile_X14Y11_FAB2RAM_D3_O0(FAB2RAM_D_O[60]),
    .Tile_X14Y11_FAB2RAM_D3_O1(FAB2RAM_D_O[61]),
    .Tile_X14Y11_FAB2RAM_D3_O2(FAB2RAM_D_O[62]),
    .Tile_X14Y11_FAB2RAM_D3_O3(FAB2RAM_D_O[63]),
    .Tile_X14Y10_FAB2RAM_D0_O0(FAB2RAM_D_O[64]),
    .Tile_X14Y10_FAB2RAM_D0_O1(FAB2RAM_D_O[65]),
    .Tile_X14Y10_FAB2RAM_D0_O2(FAB2RAM_D_O[66]),
    .Tile_X14Y10_FAB2RAM_D0_O3(FAB2RAM_D_O[67]),
    .Tile_X14Y10_FAB2RAM_D1_O0(FAB2RAM_D_O[68]),
    .Tile_X14Y10_FAB2RAM_D1_O1(FAB2RAM_D_O[69]),
    .Tile_X14Y10_FAB2RAM_D1_O2(FAB2RAM_D_O[70]),
    .Tile_X14Y10_FAB2RAM_D1_O3(FAB2RAM_D_O[71]),
    .Tile_X14Y10_FAB2RAM_D2_O0(FAB2RAM_D_O[72]),
    .Tile_X14Y10_FAB2RAM_D2_O1(FAB2RAM_D_O[73]),
    .Tile_X14Y10_FAB2RAM_D2_O2(FAB2RAM_D_O[74]),
    .Tile_X14Y10_FAB2RAM_D2_O3(FAB2RAM_D_O[75]),
    .Tile_X14Y10_FAB2RAM_D3_O0(FAB2RAM_D_O[76]),
    .Tile_X14Y10_FAB2RAM_D3_O1(FAB2RAM_D_O[77]),
    .Tile_X14Y10_FAB2RAM_D3_O2(FAB2RAM_D_O[78]),
    .Tile_X14Y10_FAB2RAM_D3_O3(FAB2RAM_D_O[79]),
    .Tile_X0Y14_B_I_top(I_top[0]),
    .Tile_X0Y14_A_I_top(I_top[1]),
    .Tile_X0Y13_B_I_top(I_top[2]),
    .Tile_X0Y13_A_I_top(I_top[3]),
    .Tile_X0Y12_B_I_top(I_top[4]),
    .Tile_X0Y12_A_I_top(I_top[5]),
    .Tile_X0Y11_B_I_top(I_top[6]),
    .Tile_X0Y11_A_I_top(I_top[7]),
    .Tile_X0Y10_B_I_top(I_top[8]),
    .Tile_X0Y10_A_I_top(I_top[9]),
    .Tile_X3Y9_OPA_I0(OPA_I[0]),
    .Tile_X3Y9_OPA_I1(OPA_I[1]),
    .Tile_X3Y9_OPA_I2(OPA_I[2]),
    .Tile_X3Y9_OPA_I3(OPA_I[3]),
    .Tile_X11Y9_OPA_I0(OPA_I[4]),
    .Tile_X11Y9_OPA_I1(OPA_I[5]),
    .Tile_X11Y9_OPA_I2(OPA_I[6]),
    .Tile_X11Y9_OPA_I3(OPA_I[7]),
    .Tile_X3Y8_OPA_I0(OPA_I[8]),
    .Tile_X3Y8_OPA_I1(OPA_I[9]),
    .Tile_X3Y8_OPA_I2(OPA_I[10]),
    .Tile_X3Y8_OPA_I3(OPA_I[11]),
    .Tile_X11Y8_OPA_I0(OPA_I[12]),
    .Tile_X11Y8_OPA_I1(OPA_I[13]),
    .Tile_X11Y8_OPA_I2(OPA_I[14]),
    .Tile_X11Y8_OPA_I3(OPA_I[15]),
    .Tile_X3Y7_OPA_I0(OPA_I[16]),
    .Tile_X3Y7_OPA_I1(OPA_I[17]),
    .Tile_X3Y7_OPA_I2(OPA_I[18]),
    .Tile_X3Y7_OPA_I3(OPA_I[19]),
    .Tile_X11Y7_OPA_I0(OPA_I[20]),
    .Tile_X11Y7_OPA_I1(OPA_I[21]),
    .Tile_X11Y7_OPA_I2(OPA_I[22]),
    .Tile_X11Y7_OPA_I3(OPA_I[23]),
    .Tile_X3Y6_OPA_I0(OPA_I[24]),
    .Tile_X3Y6_OPA_I1(OPA_I[25]),
    .Tile_X3Y6_OPA_I2(OPA_I[26]),
    .Tile_X3Y6_OPA_I3(OPA_I[27]),
    .Tile_X11Y6_OPA_I0(OPA_I[28]),
    .Tile_X11Y6_OPA_I1(OPA_I[29]),
    .Tile_X11Y6_OPA_I2(OPA_I[30]),
    .Tile_X11Y6_OPA_I3(OPA_I[31]),
    .Tile_X3Y5_OPA_I0(OPA_I[32]),
    .Tile_X3Y5_OPA_I1(OPA_I[33]),
    .Tile_X3Y5_OPA_I2(OPA_I[34]),
    .Tile_X3Y5_OPA_I3(OPA_I[35]),
    .Tile_X11Y5_OPA_I0(OPA_I[36]),
    .Tile_X11Y5_OPA_I1(OPA_I[37]),
    .Tile_X11Y5_OPA_I2(OPA_I[38]),
    .Tile_X11Y5_OPA_I3(OPA_I[39]),
    .Tile_X3Y4_OPA_I0(OPA_I[40]),
    .Tile_X3Y4_OPA_I1(OPA_I[41]),
    .Tile_X3Y4_OPA_I2(OPA_I[42]),
    .Tile_X3Y4_OPA_I3(OPA_I[43]),
    .Tile_X11Y4_OPA_I0(OPA_I[44]),
    .Tile_X11Y4_OPA_I1(OPA_I[45]),
    .Tile_X11Y4_OPA_I2(OPA_I[46]),
    .Tile_X11Y4_OPA_I3(OPA_I[47]),
    .Tile_X3Y3_OPA_I0(OPA_I[48]),
    .Tile_X3Y3_OPA_I1(OPA_I[49]),
    .Tile_X3Y3_OPA_I2(OPA_I[50]),
    .Tile_X3Y3_OPA_I3(OPA_I[51]),
    .Tile_X11Y3_OPA_I0(OPA_I[52]),
    .Tile_X11Y3_OPA_I1(OPA_I[53]),
    .Tile_X11Y3_OPA_I2(OPA_I[54]),
    .Tile_X11Y3_OPA_I3(OPA_I[55]),
    .Tile_X3Y2_OPA_I0(OPA_I[56]),
    .Tile_X3Y2_OPA_I1(OPA_I[57]),
    .Tile_X3Y2_OPA_I2(OPA_I[58]),
    .Tile_X3Y2_OPA_I3(OPA_I[59]),
    .Tile_X11Y2_OPA_I0(OPA_I[60]),
    .Tile_X11Y2_OPA_I1(OPA_I[61]),
    .Tile_X11Y2_OPA_I2(OPA_I[62]),
    .Tile_X11Y2_OPA_I3(OPA_I[63]),
    .Tile_X3Y1_OPA_I0(OPA_I[64]),
    .Tile_X3Y1_OPA_I1(OPA_I[65]),
    .Tile_X3Y1_OPA_I2(OPA_I[66]),
    .Tile_X3Y1_OPA_I3(OPA_I[67]),
    .Tile_X11Y1_OPA_I0(OPA_I[68]),
    .Tile_X11Y1_OPA_I1(OPA_I[69]),
    .Tile_X11Y1_OPA_I2(OPA_I[70]),
    .Tile_X11Y1_OPA_I3(OPA_I[71]),
    .Tile_X3Y9_OPB_I0(OPB_I[0]),
    .Tile_X3Y9_OPB_I1(OPB_I[1]),
    .Tile_X3Y9_OPB_I2(OPB_I[2]),
    .Tile_X3Y9_OPB_I3(OPB_I[3]),
    .Tile_X11Y9_OPB_I0(OPB_I[4]),
    .Tile_X11Y9_OPB_I1(OPB_I[5]),
    .Tile_X11Y9_OPB_I2(OPB_I[6]),
    .Tile_X11Y9_OPB_I3(OPB_I[7]),
    .Tile_X3Y8_OPB_I0(OPB_I[8]),
    .Tile_X3Y8_OPB_I1(OPB_I[9]),
    .Tile_X3Y8_OPB_I2(OPB_I[10]),
    .Tile_X3Y8_OPB_I3(OPB_I[11]),
    .Tile_X11Y8_OPB_I0(OPB_I[12]),
    .Tile_X11Y8_OPB_I1(OPB_I[13]),
    .Tile_X11Y8_OPB_I2(OPB_I[14]),
    .Tile_X11Y8_OPB_I3(OPB_I[15]),
    .Tile_X3Y7_OPB_I0(OPB_I[16]),
    .Tile_X3Y7_OPB_I1(OPB_I[17]),
    .Tile_X3Y7_OPB_I2(OPB_I[18]),
    .Tile_X3Y7_OPB_I3(OPB_I[19]),
    .Tile_X11Y7_OPB_I0(OPB_I[20]),
    .Tile_X11Y7_OPB_I1(OPB_I[21]),
    .Tile_X11Y7_OPB_I2(OPB_I[22]),
    .Tile_X11Y7_OPB_I3(OPB_I[23]),
    .Tile_X3Y6_OPB_I0(OPB_I[24]),
    .Tile_X3Y6_OPB_I1(OPB_I[25]),
    .Tile_X3Y6_OPB_I2(OPB_I[26]),
    .Tile_X3Y6_OPB_I3(OPB_I[27]),
    .Tile_X11Y6_OPB_I0(OPB_I[28]),
    .Tile_X11Y6_OPB_I1(OPB_I[29]),
    .Tile_X11Y6_OPB_I2(OPB_I[30]),
    .Tile_X11Y6_OPB_I3(OPB_I[31]),
    .Tile_X3Y5_OPB_I0(OPB_I[32]),
    .Tile_X3Y5_OPB_I1(OPB_I[33]),
    .Tile_X3Y5_OPB_I2(OPB_I[34]),
    .Tile_X3Y5_OPB_I3(OPB_I[35]),
    .Tile_X11Y5_OPB_I0(OPB_I[36]),
    .Tile_X11Y5_OPB_I1(OPB_I[37]),
    .Tile_X11Y5_OPB_I2(OPB_I[38]),
    .Tile_X11Y5_OPB_I3(OPB_I[39]),
    .Tile_X3Y4_OPB_I0(OPB_I[40]),
    .Tile_X3Y4_OPB_I1(OPB_I[41]),
    .Tile_X3Y4_OPB_I2(OPB_I[42]),
    .Tile_X3Y4_OPB_I3(OPB_I[43]),
    .Tile_X11Y4_OPB_I0(OPB_I[44]),
    .Tile_X11Y4_OPB_I1(OPB_I[45]),
    .Tile_X11Y4_OPB_I2(OPB_I[46]),
    .Tile_X11Y4_OPB_I3(OPB_I[47]),
    .Tile_X3Y3_OPB_I0(OPB_I[48]),
    .Tile_X3Y3_OPB_I1(OPB_I[49]),
    .Tile_X3Y3_OPB_I2(OPB_I[50]),
    .Tile_X3Y3_OPB_I3(OPB_I[51]),
    .Tile_X11Y3_OPB_I0(OPB_I[52]),
    .Tile_X11Y3_OPB_I1(OPB_I[53]),
    .Tile_X11Y3_OPB_I2(OPB_I[54]),
    .Tile_X11Y3_OPB_I3(OPB_I[55]),
    .Tile_X3Y2_OPB_I0(OPB_I[56]),
    .Tile_X3Y2_OPB_I1(OPB_I[57]),
    .Tile_X3Y2_OPB_I2(OPB_I[58]),
    .Tile_X3Y2_OPB_I3(OPB_I[59]),
    .Tile_X11Y2_OPB_I0(OPB_I[60]),
    .Tile_X11Y2_OPB_I1(OPB_I[61]),
    .Tile_X11Y2_OPB_I2(OPB_I[62]),
    .Tile_X11Y2_OPB_I3(OPB_I[63]),
    .Tile_X3Y1_OPB_I0(OPB_I[64]),
    .Tile_X3Y1_OPB_I1(OPB_I[65]),
    .Tile_X3Y1_OPB_I2(OPB_I[66]),
    .Tile_X3Y1_OPB_I3(OPB_I[67]),
    .Tile_X11Y1_OPB_I0(OPB_I[68]),
    .Tile_X11Y1_OPB_I1(OPB_I[69]),
    .Tile_X11Y1_OPB_I2(OPB_I[70]),
    .Tile_X11Y1_OPB_I3(OPB_I[71]),
    .Tile_X0Y14_B_O_top(O_top[0]),
    .Tile_X0Y14_A_O_top(O_top[1]),
    .Tile_X0Y13_B_O_top(O_top[2]),
    .Tile_X0Y13_A_O_top(O_top[3]),
    .Tile_X0Y12_B_O_top(O_top[4]),
    .Tile_X0Y12_A_O_top(O_top[5]),
    .Tile_X0Y11_B_O_top(O_top[6]),
    .Tile_X0Y11_A_O_top(O_top[7]),
    .Tile_X0Y10_B_O_top(O_top[8]),
    .Tile_X0Y10_A_O_top(O_top[9]),
    .Tile_X14Y14_RAM2FAB_D0_I0(RAM2FAB_D_I[0]),
    .Tile_X14Y14_RAM2FAB_D0_I1(RAM2FAB_D_I[1]),
    .Tile_X14Y14_RAM2FAB_D0_I2(RAM2FAB_D_I[2]),
    .Tile_X14Y14_RAM2FAB_D0_I3(RAM2FAB_D_I[3]),
    .Tile_X14Y14_RAM2FAB_D1_I0(RAM2FAB_D_I[4]),
    .Tile_X14Y14_RAM2FAB_D1_I1(RAM2FAB_D_I[5]),
    .Tile_X14Y14_RAM2FAB_D1_I2(RAM2FAB_D_I[6]),
    .Tile_X14Y14_RAM2FAB_D1_I3(RAM2FAB_D_I[7]),
    .Tile_X14Y14_RAM2FAB_D2_I0(RAM2FAB_D_I[8]),
    .Tile_X14Y14_RAM2FAB_D2_I1(RAM2FAB_D_I[9]),
    .Tile_X14Y14_RAM2FAB_D2_I2(RAM2FAB_D_I[10]),
    .Tile_X14Y14_RAM2FAB_D2_I3(RAM2FAB_D_I[11]),
    .Tile_X14Y14_RAM2FAB_D3_I0(RAM2FAB_D_I[12]),
    .Tile_X14Y14_RAM2FAB_D3_I1(RAM2FAB_D_I[13]),
    .Tile_X14Y14_RAM2FAB_D3_I2(RAM2FAB_D_I[14]),
    .Tile_X14Y14_RAM2FAB_D3_I3(RAM2FAB_D_I[15]),
    .Tile_X14Y13_RAM2FAB_D0_I0(RAM2FAB_D_I[16]),
    .Tile_X14Y13_RAM2FAB_D0_I1(RAM2FAB_D_I[17]),
    .Tile_X14Y13_RAM2FAB_D0_I2(RAM2FAB_D_I[18]),
    .Tile_X14Y13_RAM2FAB_D0_I3(RAM2FAB_D_I[19]),
    .Tile_X14Y13_RAM2FAB_D1_I0(RAM2FAB_D_I[20]),
    .Tile_X14Y13_RAM2FAB_D1_I1(RAM2FAB_D_I[21]),
    .Tile_X14Y13_RAM2FAB_D1_I2(RAM2FAB_D_I[22]),
    .Tile_X14Y13_RAM2FAB_D1_I3(RAM2FAB_D_I[23]),
    .Tile_X14Y13_RAM2FAB_D2_I0(RAM2FAB_D_I[24]),
    .Tile_X14Y13_RAM2FAB_D2_I1(RAM2FAB_D_I[25]),
    .Tile_X14Y13_RAM2FAB_D2_I2(RAM2FAB_D_I[26]),
    .Tile_X14Y13_RAM2FAB_D2_I3(RAM2FAB_D_I[27]),
    .Tile_X14Y13_RAM2FAB_D3_I0(RAM2FAB_D_I[28]),
    .Tile_X14Y13_RAM2FAB_D3_I1(RAM2FAB_D_I[29]),
    .Tile_X14Y13_RAM2FAB_D3_I2(RAM2FAB_D_I[30]),
    .Tile_X14Y13_RAM2FAB_D3_I3(RAM2FAB_D_I[31]),
    .Tile_X14Y12_RAM2FAB_D0_I0(RAM2FAB_D_I[32]),
    .Tile_X14Y12_RAM2FAB_D0_I1(RAM2FAB_D_I[33]),
    .Tile_X14Y12_RAM2FAB_D0_I2(RAM2FAB_D_I[34]),
    .Tile_X14Y12_RAM2FAB_D0_I3(RAM2FAB_D_I[35]),
    .Tile_X14Y12_RAM2FAB_D1_I0(RAM2FAB_D_I[36]),
    .Tile_X14Y12_RAM2FAB_D1_I1(RAM2FAB_D_I[37]),
    .Tile_X14Y12_RAM2FAB_D1_I2(RAM2FAB_D_I[38]),
    .Tile_X14Y12_RAM2FAB_D1_I3(RAM2FAB_D_I[39]),
    .Tile_X14Y12_RAM2FAB_D2_I0(RAM2FAB_D_I[40]),
    .Tile_X14Y12_RAM2FAB_D2_I1(RAM2FAB_D_I[41]),
    .Tile_X14Y12_RAM2FAB_D2_I2(RAM2FAB_D_I[42]),
    .Tile_X14Y12_RAM2FAB_D2_I3(RAM2FAB_D_I[43]),
    .Tile_X14Y12_RAM2FAB_D3_I0(RAM2FAB_D_I[44]),
    .Tile_X14Y12_RAM2FAB_D3_I1(RAM2FAB_D_I[45]),
    .Tile_X14Y12_RAM2FAB_D3_I2(RAM2FAB_D_I[46]),
    .Tile_X14Y12_RAM2FAB_D3_I3(RAM2FAB_D_I[47]),
    .Tile_X14Y11_RAM2FAB_D0_I0(RAM2FAB_D_I[48]),
    .Tile_X14Y11_RAM2FAB_D0_I1(RAM2FAB_D_I[49]),
    .Tile_X14Y11_RAM2FAB_D0_I2(RAM2FAB_D_I[50]),
    .Tile_X14Y11_RAM2FAB_D0_I3(RAM2FAB_D_I[51]),
    .Tile_X14Y11_RAM2FAB_D1_I0(RAM2FAB_D_I[52]),
    .Tile_X14Y11_RAM2FAB_D1_I1(RAM2FAB_D_I[53]),
    .Tile_X14Y11_RAM2FAB_D1_I2(RAM2FAB_D_I[54]),
    .Tile_X14Y11_RAM2FAB_D1_I3(RAM2FAB_D_I[55]),
    .Tile_X14Y11_RAM2FAB_D2_I0(RAM2FAB_D_I[56]),
    .Tile_X14Y11_RAM2FAB_D2_I1(RAM2FAB_D_I[57]),
    .Tile_X14Y11_RAM2FAB_D2_I2(RAM2FAB_D_I[58]),
    .Tile_X14Y11_RAM2FAB_D2_I3(RAM2FAB_D_I[59]),
    .Tile_X14Y11_RAM2FAB_D3_I0(RAM2FAB_D_I[60]),
    .Tile_X14Y11_RAM2FAB_D3_I1(RAM2FAB_D_I[61]),
    .Tile_X14Y11_RAM2FAB_D3_I2(RAM2FAB_D_I[62]),
    .Tile_X14Y11_RAM2FAB_D3_I3(RAM2FAB_D_I[63]),
    .Tile_X14Y10_RAM2FAB_D0_I0(RAM2FAB_D_I[64]),
    .Tile_X14Y10_RAM2FAB_D0_I1(RAM2FAB_D_I[65]),
    .Tile_X14Y10_RAM2FAB_D0_I2(RAM2FAB_D_I[66]),
    .Tile_X14Y10_RAM2FAB_D0_I3(RAM2FAB_D_I[67]),
    .Tile_X14Y10_RAM2FAB_D1_I0(RAM2FAB_D_I[68]),
    .Tile_X14Y10_RAM2FAB_D1_I1(RAM2FAB_D_I[69]),
    .Tile_X14Y10_RAM2FAB_D1_I2(RAM2FAB_D_I[70]),
    .Tile_X14Y10_RAM2FAB_D1_I3(RAM2FAB_D_I[71]),
    .Tile_X14Y10_RAM2FAB_D2_I0(RAM2FAB_D_I[72]),
    .Tile_X14Y10_RAM2FAB_D2_I1(RAM2FAB_D_I[73]),
    .Tile_X14Y10_RAM2FAB_D2_I2(RAM2FAB_D_I[74]),
    .Tile_X14Y10_RAM2FAB_D2_I3(RAM2FAB_D_I[75]),
    .Tile_X14Y10_RAM2FAB_D3_I0(RAM2FAB_D_I[76]),
    .Tile_X14Y10_RAM2FAB_D3_I1(RAM2FAB_D_I[77]),
    .Tile_X14Y10_RAM2FAB_D3_I2(RAM2FAB_D_I[78]),
    .Tile_X14Y10_RAM2FAB_D3_I3(RAM2FAB_D_I[79]),
    .Tile_X3Y9_RES0_O0(RES0_O[0]),
    .Tile_X3Y9_RES0_O1(RES0_O[1]),
    .Tile_X3Y9_RES0_O2(RES0_O[2]),
    .Tile_X3Y9_RES0_O3(RES0_O[3]),
    .Tile_X11Y9_RES0_O0(RES0_O[4]),
    .Tile_X11Y9_RES0_O1(RES0_O[5]),
    .Tile_X11Y9_RES0_O2(RES0_O[6]),
    .Tile_X11Y9_RES0_O3(RES0_O[7]),
    .Tile_X3Y8_RES0_O0(RES0_O[8]),
    .Tile_X3Y8_RES0_O1(RES0_O[9]),
    .Tile_X3Y8_RES0_O2(RES0_O[10]),
    .Tile_X3Y8_RES0_O3(RES0_O[11]),
    .Tile_X11Y8_RES0_O0(RES0_O[12]),
    .Tile_X11Y8_RES0_O1(RES0_O[13]),
    .Tile_X11Y8_RES0_O2(RES0_O[14]),
    .Tile_X11Y8_RES0_O3(RES0_O[15]),
    .Tile_X3Y7_RES0_O0(RES0_O[16]),
    .Tile_X3Y7_RES0_O1(RES0_O[17]),
    .Tile_X3Y7_RES0_O2(RES0_O[18]),
    .Tile_X3Y7_RES0_O3(RES0_O[19]),
    .Tile_X11Y7_RES0_O0(RES0_O[20]),
    .Tile_X11Y7_RES0_O1(RES0_O[21]),
    .Tile_X11Y7_RES0_O2(RES0_O[22]),
    .Tile_X11Y7_RES0_O3(RES0_O[23]),
    .Tile_X3Y6_RES0_O0(RES0_O[24]),
    .Tile_X3Y6_RES0_O1(RES0_O[25]),
    .Tile_X3Y6_RES0_O2(RES0_O[26]),
    .Tile_X3Y6_RES0_O3(RES0_O[27]),
    .Tile_X11Y6_RES0_O0(RES0_O[28]),
    .Tile_X11Y6_RES0_O1(RES0_O[29]),
    .Tile_X11Y6_RES0_O2(RES0_O[30]),
    .Tile_X11Y6_RES0_O3(RES0_O[31]),
    .Tile_X3Y5_RES0_O0(RES0_O[32]),
    .Tile_X3Y5_RES0_O1(RES0_O[33]),
    .Tile_X3Y5_RES0_O2(RES0_O[34]),
    .Tile_X3Y5_RES0_O3(RES0_O[35]),
    .Tile_X11Y5_RES0_O0(RES0_O[36]),
    .Tile_X11Y5_RES0_O1(RES0_O[37]),
    .Tile_X11Y5_RES0_O2(RES0_O[38]),
    .Tile_X11Y5_RES0_O3(RES0_O[39]),
    .Tile_X3Y4_RES0_O0(RES0_O[40]),
    .Tile_X3Y4_RES0_O1(RES0_O[41]),
    .Tile_X3Y4_RES0_O2(RES0_O[42]),
    .Tile_X3Y4_RES0_O3(RES0_O[43]),
    .Tile_X11Y4_RES0_O0(RES0_O[44]),
    .Tile_X11Y4_RES0_O1(RES0_O[45]),
    .Tile_X11Y4_RES0_O2(RES0_O[46]),
    .Tile_X11Y4_RES0_O3(RES0_O[47]),
    .Tile_X3Y3_RES0_O0(RES0_O[48]),
    .Tile_X3Y3_RES0_O1(RES0_O[49]),
    .Tile_X3Y3_RES0_O2(RES0_O[50]),
    .Tile_X3Y3_RES0_O3(RES0_O[51]),
    .Tile_X11Y3_RES0_O0(RES0_O[52]),
    .Tile_X11Y3_RES0_O1(RES0_O[53]),
    .Tile_X11Y3_RES0_O2(RES0_O[54]),
    .Tile_X11Y3_RES0_O3(RES0_O[55]),
    .Tile_X3Y2_RES0_O0(RES0_O[56]),
    .Tile_X3Y2_RES0_O1(RES0_O[57]),
    .Tile_X3Y2_RES0_O2(RES0_O[58]),
    .Tile_X3Y2_RES0_O3(RES0_O[59]),
    .Tile_X11Y2_RES0_O0(RES0_O[60]),
    .Tile_X11Y2_RES0_O1(RES0_O[61]),
    .Tile_X11Y2_RES0_O2(RES0_O[62]),
    .Tile_X11Y2_RES0_O3(RES0_O[63]),
    .Tile_X3Y1_RES0_O0(RES0_O[64]),
    .Tile_X3Y1_RES0_O1(RES0_O[65]),
    .Tile_X3Y1_RES0_O2(RES0_O[66]),
    .Tile_X3Y1_RES0_O3(RES0_O[67]),
    .Tile_X11Y1_RES0_O0(RES0_O[68]),
    .Tile_X11Y1_RES0_O1(RES0_O[69]),
    .Tile_X11Y1_RES0_O2(RES0_O[70]),
    .Tile_X11Y1_RES0_O3(RES0_O[71]),
    .Tile_X3Y9_RES1_O0(RES1_O[0]),
    .Tile_X3Y9_RES1_O1(RES1_O[1]),
    .Tile_X3Y9_RES1_O2(RES1_O[2]),
    .Tile_X3Y9_RES1_O3(RES1_O[3]),
    .Tile_X11Y9_RES1_O0(RES1_O[4]),
    .Tile_X11Y9_RES1_O1(RES1_O[5]),
    .Tile_X11Y9_RES1_O2(RES1_O[6]),
    .Tile_X11Y9_RES1_O3(RES1_O[7]),
    .Tile_X3Y8_RES1_O0(RES1_O[8]),
    .Tile_X3Y8_RES1_O1(RES1_O[9]),
    .Tile_X3Y8_RES1_O2(RES1_O[10]),
    .Tile_X3Y8_RES1_O3(RES1_O[11]),
    .Tile_X11Y8_RES1_O0(RES1_O[12]),
    .Tile_X11Y8_RES1_O1(RES1_O[13]),
    .Tile_X11Y8_RES1_O2(RES1_O[14]),
    .Tile_X11Y8_RES1_O3(RES1_O[15]),
    .Tile_X3Y7_RES1_O0(RES1_O[16]),
    .Tile_X3Y7_RES1_O1(RES1_O[17]),
    .Tile_X3Y7_RES1_O2(RES1_O[18]),
    .Tile_X3Y7_RES1_O3(RES1_O[19]),
    .Tile_X11Y7_RES1_O0(RES1_O[20]),
    .Tile_X11Y7_RES1_O1(RES1_O[21]),
    .Tile_X11Y7_RES1_O2(RES1_O[22]),
    .Tile_X11Y7_RES1_O3(RES1_O[23]),
    .Tile_X3Y6_RES1_O0(RES1_O[24]),
    .Tile_X3Y6_RES1_O1(RES1_O[25]),
    .Tile_X3Y6_RES1_O2(RES1_O[26]),
    .Tile_X3Y6_RES1_O3(RES1_O[27]),
    .Tile_X11Y6_RES1_O0(RES1_O[28]),
    .Tile_X11Y6_RES1_O1(RES1_O[29]),
    .Tile_X11Y6_RES1_O2(RES1_O[30]),
    .Tile_X11Y6_RES1_O3(RES1_O[31]),
    .Tile_X3Y5_RES1_O0(RES1_O[32]),
    .Tile_X3Y5_RES1_O1(RES1_O[33]),
    .Tile_X3Y5_RES1_O2(RES1_O[34]),
    .Tile_X3Y5_RES1_O3(RES1_O[35]),
    .Tile_X11Y5_RES1_O0(RES1_O[36]),
    .Tile_X11Y5_RES1_O1(RES1_O[37]),
    .Tile_X11Y5_RES1_O2(RES1_O[38]),
    .Tile_X11Y5_RES1_O3(RES1_O[39]),
    .Tile_X3Y4_RES1_O0(RES1_O[40]),
    .Tile_X3Y4_RES1_O1(RES1_O[41]),
    .Tile_X3Y4_RES1_O2(RES1_O[42]),
    .Tile_X3Y4_RES1_O3(RES1_O[43]),
    .Tile_X11Y4_RES1_O0(RES1_O[44]),
    .Tile_X11Y4_RES1_O1(RES1_O[45]),
    .Tile_X11Y4_RES1_O2(RES1_O[46]),
    .Tile_X11Y4_RES1_O3(RES1_O[47]),
    .Tile_X3Y3_RES1_O0(RES1_O[48]),
    .Tile_X3Y3_RES1_O1(RES1_O[49]),
    .Tile_X3Y3_RES1_O2(RES1_O[50]),
    .Tile_X3Y3_RES1_O3(RES1_O[51]),
    .Tile_X11Y3_RES1_O0(RES1_O[52]),
    .Tile_X11Y3_RES1_O1(RES1_O[53]),
    .Tile_X11Y3_RES1_O2(RES1_O[54]),
    .Tile_X11Y3_RES1_O3(RES1_O[55]),
    .Tile_X3Y2_RES1_O0(RES1_O[56]),
    .Tile_X3Y2_RES1_O1(RES1_O[57]),
    .Tile_X3Y2_RES1_O2(RES1_O[58]),
    .Tile_X3Y2_RES1_O3(RES1_O[59]),
    .Tile_X11Y2_RES1_O0(RES1_O[60]),
    .Tile_X11Y2_RES1_O1(RES1_O[61]),
    .Tile_X11Y2_RES1_O2(RES1_O[62]),
    .Tile_X11Y2_RES1_O3(RES1_O[63]),
    .Tile_X3Y1_RES1_O0(RES1_O[64]),
    .Tile_X3Y1_RES1_O1(RES1_O[65]),
    .Tile_X3Y1_RES1_O2(RES1_O[66]),
    .Tile_X3Y1_RES1_O3(RES1_O[67]),
    .Tile_X11Y1_RES1_O0(RES1_O[68]),
    .Tile_X11Y1_RES1_O1(RES1_O[69]),
    .Tile_X11Y1_RES1_O2(RES1_O[70]),
    .Tile_X11Y1_RES1_O3(RES1_O[71]),
    .Tile_X3Y9_RES2_O0(RES2_O[0]),
    .Tile_X3Y9_RES2_O1(RES2_O[1]),
    .Tile_X3Y9_RES2_O2(RES2_O[2]),
    .Tile_X3Y9_RES2_O3(RES2_O[3]),
    .Tile_X11Y9_RES2_O0(RES2_O[4]),
    .Tile_X11Y9_RES2_O1(RES2_O[5]),
    .Tile_X11Y9_RES2_O2(RES2_O[6]),
    .Tile_X11Y9_RES2_O3(RES2_O[7]),
    .Tile_X3Y8_RES2_O0(RES2_O[8]),
    .Tile_X3Y8_RES2_O1(RES2_O[9]),
    .Tile_X3Y8_RES2_O2(RES2_O[10]),
    .Tile_X3Y8_RES2_O3(RES2_O[11]),
    .Tile_X11Y8_RES2_O0(RES2_O[12]),
    .Tile_X11Y8_RES2_O1(RES2_O[13]),
    .Tile_X11Y8_RES2_O2(RES2_O[14]),
    .Tile_X11Y8_RES2_O3(RES2_O[15]),
    .Tile_X3Y7_RES2_O0(RES2_O[16]),
    .Tile_X3Y7_RES2_O1(RES2_O[17]),
    .Tile_X3Y7_RES2_O2(RES2_O[18]),
    .Tile_X3Y7_RES2_O3(RES2_O[19]),
    .Tile_X11Y7_RES2_O0(RES2_O[20]),
    .Tile_X11Y7_RES2_O1(RES2_O[21]),
    .Tile_X11Y7_RES2_O2(RES2_O[22]),
    .Tile_X11Y7_RES2_O3(RES2_O[23]),
    .Tile_X3Y6_RES2_O0(RES2_O[24]),
    .Tile_X3Y6_RES2_O1(RES2_O[25]),
    .Tile_X3Y6_RES2_O2(RES2_O[26]),
    .Tile_X3Y6_RES2_O3(RES2_O[27]),
    .Tile_X11Y6_RES2_O0(RES2_O[28]),
    .Tile_X11Y6_RES2_O1(RES2_O[29]),
    .Tile_X11Y6_RES2_O2(RES2_O[30]),
    .Tile_X11Y6_RES2_O3(RES2_O[31]),
    .Tile_X3Y5_RES2_O0(RES2_O[32]),
    .Tile_X3Y5_RES2_O1(RES2_O[33]),
    .Tile_X3Y5_RES2_O2(RES2_O[34]),
    .Tile_X3Y5_RES2_O3(RES2_O[35]),
    .Tile_X11Y5_RES2_O0(RES2_O[36]),
    .Tile_X11Y5_RES2_O1(RES2_O[37]),
    .Tile_X11Y5_RES2_O2(RES2_O[38]),
    .Tile_X11Y5_RES2_O3(RES2_O[39]),
    .Tile_X3Y4_RES2_O0(RES2_O[40]),
    .Tile_X3Y4_RES2_O1(RES2_O[41]),
    .Tile_X3Y4_RES2_O2(RES2_O[42]),
    .Tile_X3Y4_RES2_O3(RES2_O[43]),
    .Tile_X11Y4_RES2_O0(RES2_O[44]),
    .Tile_X11Y4_RES2_O1(RES2_O[45]),
    .Tile_X11Y4_RES2_O2(RES2_O[46]),
    .Tile_X11Y4_RES2_O3(RES2_O[47]),
    .Tile_X3Y3_RES2_O0(RES2_O[48]),
    .Tile_X3Y3_RES2_O1(RES2_O[49]),
    .Tile_X3Y3_RES2_O2(RES2_O[50]),
    .Tile_X3Y3_RES2_O3(RES2_O[51]),
    .Tile_X11Y3_RES2_O0(RES2_O[52]),
    .Tile_X11Y3_RES2_O1(RES2_O[53]),
    .Tile_X11Y3_RES2_O2(RES2_O[54]),
    .Tile_X11Y3_RES2_O3(RES2_O[55]),
    .Tile_X3Y2_RES2_O0(RES2_O[56]),
    .Tile_X3Y2_RES2_O1(RES2_O[57]),
    .Tile_X3Y2_RES2_O2(RES2_O[58]),
    .Tile_X3Y2_RES2_O3(RES2_O[59]),
    .Tile_X11Y2_RES2_O0(RES2_O[60]),
    .Tile_X11Y2_RES2_O1(RES2_O[61]),
    .Tile_X11Y2_RES2_O2(RES2_O[62]),
    .Tile_X11Y2_RES2_O3(RES2_O[63]),
    .Tile_X3Y1_RES2_O0(RES2_O[64]),
    .Tile_X3Y1_RES2_O1(RES2_O[65]),
    .Tile_X3Y1_RES2_O2(RES2_O[66]),
    .Tile_X3Y1_RES2_O3(RES2_O[67]),
    .Tile_X11Y1_RES2_O0(RES2_O[68]),
    .Tile_X11Y1_RES2_O1(RES2_O[69]),
    .Tile_X11Y1_RES2_O2(RES2_O[70]),
    .Tile_X11Y1_RES2_O3(RES2_O[71]),
    .Tile_X0Y14_B_T_top(T_top[0]),
    .Tile_X0Y14_A_T_top(T_top[1]),
    .Tile_X0Y13_B_T_top(T_top[2]),
    .Tile_X0Y13_A_T_top(T_top[3]),
    .Tile_X0Y12_B_T_top(T_top[4]),
    .Tile_X0Y12_A_T_top(T_top[5]),
    .Tile_X0Y11_B_T_top(T_top[6]),
    .Tile_X0Y11_A_T_top(T_top[7]),
    .Tile_X0Y10_B_T_top(T_top[8]),
    .Tile_X0Y10_A_T_top(T_top[9]),
    .UserCLK(CLK),
    .FrameData(FrameData),
    .FrameStrobe(FrameSelect)
);*/


// BlockRAM_1KB Inst_BlockRAM_0 (
//     .clk(CLK),
//     .rd_addr(FAB2RAM_A_O[7:0]),
//     .rd_data(RAM2FAB_D_I[31:0]),
//     .wr_addr(FAB2RAM_A_O[15:8]),
//     .wr_data(FAB2RAM_D_O[31:0]),
//     .C0(FAB2RAM_C_O[0]),
//     .C1(FAB2RAM_C_O[1]),
//     .C2(FAB2RAM_C_O[2]),
//     .C3(FAB2RAM_C_O[3]),
//     .C4(FAB2RAM_C_O[4]),
//     .C5(FAB2RAM_C_O[5])
// );

// BlockRAM_1KB Inst_BlockRAM_1 (
//     .clk(CLK),
//     .rd_addr(FAB2RAM_A_O[23:16]),
//     .rd_data(RAM2FAB_D_I[63:32]),
//     .wr_addr(FAB2RAM_A_O[31:24]),
//     .wr_data(FAB2RAM_D_O[63:32]),
//     .C0(FAB2RAM_C_O[8]),
//     .C1(FAB2RAM_C_O[9]),
//     .C2(FAB2RAM_C_O[10]),
//     .C3(FAB2RAM_C_O[11]),
//     .C4(FAB2RAM_C_O[12]),
//     .C5(FAB2RAM_C_O[13])
// );

// BlockRAM_1KB Inst_BlockRAM_2 (
//     .clk(CLK),
//     .rd_addr(FAB2RAM_A_O[39:32]),
//     .rd_data(RAM2FAB_D_I[95:64]),
//     .wr_addr(FAB2RAM_A_O[47:40]),
//     .wr_data(FAB2RAM_D_O[95:64]),
//     .C0(FAB2RAM_C_O[16]),
//     .C1(FAB2RAM_C_O[17]),
//     .C2(FAB2RAM_C_O[18]),
//     .C3(FAB2RAM_C_O[19]),
//     .C4(FAB2RAM_C_O[20]),
//     .C5(FAB2RAM_C_O[21])
// );

// BlockRAM_1KB Inst_BlockRAM_3 (
//     .clk(CLK),
//     .rd_addr(FAB2RAM_A_O[55:48]),
//     .rd_data(RAM2FAB_D_I[127:96]),
//     .wr_addr(FAB2RAM_A_O[63:56]),
//     .wr_data(FAB2RAM_D_O[127:96]),
//     .C0(FAB2RAM_C_O[24]),
//     .C1(FAB2RAM_C_O[25]),
//     .C2(FAB2RAM_C_O[26]),
//     .C3(FAB2RAM_C_O[27]),
//     .C4(FAB2RAM_C_O[28]),
//     .C5(FAB2RAM_C_O[29])
// );

// BlockRAM_1KB Inst_BlockRAM_4 (
//     .clk(CLK),
//     .rd_addr(FAB2RAM_A_O[71:64]),
//     .rd_data(RAM2FAB_D_I[159:128]),
//     .wr_addr(FAB2RAM_A_O[79:72]),
//     .wr_data(FAB2RAM_D_O[159:128]),
//     .C0(FAB2RAM_C_O[32]),
//     .C1(FAB2RAM_C_O[33]),
//     .C2(FAB2RAM_C_O[34]),
//     .C3(FAB2RAM_C_O[35]),
//     .C4(FAB2RAM_C_O[36]),
//     .C5(FAB2RAM_C_O[37])
// );

// BlockRAM_1KB Inst_BlockRAM_5 (
//     .clk(CLK),
//     .rd_addr(FAB2RAM_A_O[87:80]),
//     .rd_data(RAM2FAB_D_I[191:160]),
//     .wr_addr(FAB2RAM_A_O[95:88]),
//     .wr_data(FAB2RAM_D_O[191:160]),
//     .C0(FAB2RAM_C_O[40]),
//     .C1(FAB2RAM_C_O[41]),
//     .C2(FAB2RAM_C_O[42]),
//     .C3(FAB2RAM_C_O[43]),
//     .C4(FAB2RAM_C_O[44]),
//     .C5(FAB2RAM_C_O[45])
// );

// BlockRAM_1KB Inst_BlockRAM_6 (
//     .clk(CLK),
//     .rd_addr(FAB2RAM_A_O[103:96]),
//     .rd_data(RAM2FAB_D_I[223:192]),
//     .wr_addr(FAB2RAM_A_O[111:104]),
//     .wr_data(FAB2RAM_D_O[223:192]),
//     .C0(FAB2RAM_C_O[48]),
//     .C1(FAB2RAM_C_O[49]),
//     .C2(FAB2RAM_C_O[50]),
//     .C3(FAB2RAM_C_O[51]),
//     .C4(FAB2RAM_C_O[52]),
//     .C5(FAB2RAM_C_O[53])
// );

assign FrameData = {32'h12345678,FrameRegister,32'h12345678};
endmodule