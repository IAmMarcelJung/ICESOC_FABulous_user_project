module top_wrapper;

wire clk;
(* keep *) Global_Clock clk_i (.CLK(clk));

//(* keep, BEL="X0Y14.D" *) Config_access bel_X0Y14_D ();
//(* keep, BEL="X0Y14.C" *) Config_access bel_X0Y14_C ();
(* keep, BEL="X0Y14.B" *) IO_1_bidirectional_frame_config_pass bel_X0Y14_B (.I(IO_1_bidirectional_frame_config_pass_I[0]), .T(IO_1_bidirectional_frame_config_pass_T[0]), .O(IO_1_bidirectional_frame_config_pass_O[0]), .Q(IO_1_bidirectional_frame_config_pass_Q[0]));
(* keep, BEL="X0Y14.A" *) IO_1_bidirectional_frame_config_pass bel_X0Y14_A (.I(IO_1_bidirectional_frame_config_pass_I[1]), .T(IO_1_bidirectional_frame_config_pass_T[1]), .O(IO_1_bidirectional_frame_config_pass_O[1]), .Q(IO_1_bidirectional_frame_config_pass_Q[1]));
//(* keep, BEL="X0Y13.D" *) Config_access bel_X0Y13_D ();
//(* keep, BEL="X0Y13.C" *) Config_access bel_X0Y13_C ();
(* keep, BEL="X0Y13.B" *) IO_1_bidirectional_frame_config_pass bel_X0Y13_B (.I(IO_1_bidirectional_frame_config_pass_I[2]), .T(IO_1_bidirectional_frame_config_pass_T[2]), .O(IO_1_bidirectional_frame_config_pass_O[2]), .Q(IO_1_bidirectional_frame_config_pass_Q[2]));
(* keep, BEL="X0Y13.A" *) IO_1_bidirectional_frame_config_pass bel_X0Y13_A (.I(IO_1_bidirectional_frame_config_pass_I[3]), .T(IO_1_bidirectional_frame_config_pass_T[3]), .O(IO_1_bidirectional_frame_config_pass_O[3]), .Q(IO_1_bidirectional_frame_config_pass_Q[3]));
//(* keep, BEL="X0Y12.D" *) Config_access bel_X0Y12_D ();
//(* keep, BEL="X0Y12.C" *) Config_access bel_X0Y12_C ();
(* keep, BEL="X0Y12.B" *) IO_1_bidirectional_frame_config_pass bel_X0Y12_B (.I(IO_1_bidirectional_frame_config_pass_I[4]), .T(IO_1_bidirectional_frame_config_pass_T[4]), .O(IO_1_bidirectional_frame_config_pass_O[4]), .Q(IO_1_bidirectional_frame_config_pass_Q[4]));
(* keep, BEL="X0Y12.A" *) IO_1_bidirectional_frame_config_pass bel_X0Y12_A (.I(IO_1_bidirectional_frame_config_pass_I[5]), .T(IO_1_bidirectional_frame_config_pass_T[5]), .O(IO_1_bidirectional_frame_config_pass_O[5]), .Q(IO_1_bidirectional_frame_config_pass_Q[5]));
//(* keep, BEL="X0Y11.D" *) Config_access bel_X0Y11_D ();
//(* keep, BEL="X0Y11.C" *) Config_access bel_X0Y11_C ();
(* keep, BEL="X0Y11.B" *) IO_1_bidirectional_frame_config_pass bel_X0Y11_B (.I(IO_1_bidirectional_frame_config_pass_I[6]), .T(IO_1_bidirectional_frame_config_pass_T[6]), .O(IO_1_bidirectional_frame_config_pass_O[6]), .Q(IO_1_bidirectional_frame_config_pass_Q[6]));
(* keep, BEL="X0Y11.A" *) IO_1_bidirectional_frame_config_pass bel_X0Y11_A (.I(IO_1_bidirectional_frame_config_pass_I[7]), .T(IO_1_bidirectional_frame_config_pass_T[7]), .O(IO_1_bidirectional_frame_config_pass_O[7]), .Q(IO_1_bidirectional_frame_config_pass_Q[7]));
//(* keep, BEL="X0Y10.D" *) Config_access bel_X0Y10_D ();
//(* keep, BEL="X0Y10.C" *) Config_access bel_X0Y10_C ();
(* keep, BEL="X0Y10.B" *) IO_1_bidirectional_frame_config_pass bel_X0Y10_B (.I(IO_1_bidirectional_frame_config_pass_I[8]), .T(IO_1_bidirectional_frame_config_pass_T[8]), .O(IO_1_bidirectional_frame_config_pass_O[8]), .Q(IO_1_bidirectional_frame_config_pass_Q[8]));
(* keep, BEL="X0Y10.A" *) IO_1_bidirectional_frame_config_pass bel_X0Y10_A (.I(IO_1_bidirectional_frame_config_pass_I[9]), .T(IO_1_bidirectional_frame_config_pass_T[9]), .O(IO_1_bidirectional_frame_config_pass_O[9]), .Q(IO_1_bidirectional_frame_config_pass_Q[9]));
(* keep, BEL="X3Y9.RES2" *) OutPass4_frame_config bel_X3Y9_RES2 (.I0(W_RES2[3]), .I1(W_RES2[2]), .I2(W_RES2[1]), .I3(W_RES2[0]));
(* keep, BEL="X3Y9.RES1" *) OutPass4_frame_config bel_X3Y9_RES1 (.I0(W_RES1[3]), .I1(W_RES1[2]), .I2(W_RES1[1]), .I3(W_RES1[0]));
(* keep, BEL="X3Y9.RES0" *) OutPass4_frame_config bel_X3Y9_RES0 (.I0(W_RES0[3]), .I1(W_RES0[2]), .I2(W_RES0[1]), .I3(W_RES0[0]));
(* keep, BEL="X3Y9.OPB" *) InPass4_frame_config bel_X3Y9_OPB (.O0(W_OPB[3]), .O1(W_OPB[2]), .O2(W_OPB[1]), .O3(W_OPB[0]));
(* keep, BEL="X3Y9.OPA" *) InPass4_frame_config bel_X3Y9_OPA (.O0(W_OPA[3]), .O1(W_OPA[2]), .O2(W_OPA[1]), .O3(W_OPA[0]));
(* keep, BEL="X3Y8.RES2" *) OutPass4_frame_config bel_X3Y8_RES2 (.I0(W_RES2[7]), .I1(W_RES2[6]), .I2(W_RES2[5]), .I3(W_RES2[4]));
(* keep, BEL="X3Y8.RES1" *) OutPass4_frame_config bel_X3Y8_RES1 (.I0(W_RES1[7]), .I1(W_RES1[6]), .I2(W_RES1[5]), .I3(W_RES1[4]));
(* keep, BEL="X3Y8.RES0" *) OutPass4_frame_config bel_X3Y8_RES0 (.I0(W_RES0[7]), .I1(W_RES0[6]), .I2(W_RES0[5]), .I3(W_RES0[4]));
(* keep, BEL="X3Y8.OPB" *) InPass4_frame_config bel_X3Y8_OPB (.O0(W_OPB[7]), .O1(W_OPB[6]), .O2(W_OPB[5]), .O3(W_OPB[4]));
(* keep, BEL="X3Y8.OPA" *) InPass4_frame_config bel_X3Y8_OPA (.O0(W_OPA[7]), .O1(W_OPA[6]), .O2(W_OPA[5]), .O3(W_OPA[4]));
(* keep, BEL="X3Y7.RES2" *) OutPass4_frame_config bel_X3Y7_RES2 (.I0(W_RES2[11]), .I1(W_RES2[10]), .I2(W_RES2[9]), .I3(W_RES2[8]));
(* keep, BEL="X3Y7.RES1" *) OutPass4_frame_config bel_X3Y7_RES1 (.I0(W_RES1[11]), .I1(W_RES1[10]), .I2(W_RES1[9]), .I3(W_RES1[8]));
(* keep, BEL="X3Y7.RES0" *) OutPass4_frame_config bel_X3Y7_RES0 (.I0(W_RES0[11]), .I1(W_RES0[10]), .I2(W_RES0[9]), .I3(W_RES0[8]));
(* keep, BEL="X3Y7.OPB" *) InPass4_frame_config bel_X3Y7_OPB (.O0(W_OPB[11]), .O1(W_OPB[10]), .O2(W_OPB[9]), .O3(W_OPB[8]));
(* keep, BEL="X3Y7.OPA" *) InPass4_frame_config bel_X3Y7_OPA (.O0(W_OPA[11]), .O1(W_OPA[10]), .O2(W_OPA[9]), .O3(W_OPA[8]));
(* keep, BEL="X3Y6.RES2" *) OutPass4_frame_config bel_X3Y6_RES2 (.I0(W_RES2[15]), .I1(W_RES2[14]), .I2(W_RES2[13]), .I3(W_RES2[12]));
(* keep, BEL="X3Y6.RES1" *) OutPass4_frame_config bel_X3Y6_RES1 (.I0(W_RES1[15]), .I1(W_RES1[14]), .I2(W_RES1[13]), .I3(W_RES1[12]));
(* keep, BEL="X3Y6.RES0" *) OutPass4_frame_config bel_X3Y6_RES0 (.I0(W_RES0[15]), .I1(W_RES0[14]), .I2(W_RES0[13]), .I3(W_RES0[12]));
(* keep, BEL="X3Y6.OPB" *) InPass4_frame_config bel_X3Y6_OPB (.O0(W_OPB[15]), .O1(W_OPB[14]), .O2(W_OPB[13]), .O3(W_OPB[12]));
(* keep, BEL="X3Y6.OPA" *) InPass4_frame_config bel_X3Y6_OPA (.O0(W_OPA[15]), .O1(W_OPA[14]), .O2(W_OPA[13]), .O3(W_OPA[12]));
(* keep, BEL="X3Y5.RES2" *) OutPass4_frame_config bel_X3Y5_RES2 (.I0(W_RES2[19]), .I1(W_RES2[18]), .I2(W_RES2[17]), .I3(W_RES2[16]));
(* keep, BEL="X3Y5.RES1" *) OutPass4_frame_config bel_X3Y5_RES1 (.I0(W_RES1[19]), .I1(W_RES1[18]), .I2(W_RES1[17]), .I3(W_RES1[16]));
(* keep, BEL="X3Y5.RES0" *) OutPass4_frame_config bel_X3Y5_RES0 (.I0(W_RES0[19]), .I1(W_RES0[18]), .I2(W_RES0[17]), .I3(W_RES0[16]));
(* keep, BEL="X3Y5.OPB" *) InPass4_frame_config bel_X3Y5_OPB (.O0(W_OPB[19]), .O1(W_OPB[18]), .O2(W_OPB[17]), .O3(W_OPB[16]));
(* keep, BEL="X3Y5.OPA" *) InPass4_frame_config bel_X3Y5_OPA (.O0(W_OPA[19]), .O1(W_OPA[18]), .O2(W_OPA[17]), .O3(W_OPA[16]));
(* keep, BEL="X3Y4.RES2" *) OutPass4_frame_config bel_X3Y4_RES2 (.I0(W_RES2[23]), .I1(W_RES2[22]), .I2(W_RES2[21]), .I3(W_RES2[20]));
(* keep, BEL="X3Y4.RES1" *) OutPass4_frame_config bel_X3Y4_RES1 (.I0(W_RES1[23]), .I1(W_RES1[22]), .I2(W_RES1[21]), .I3(W_RES1[20]));
(* keep, BEL="X3Y4.RES0" *) OutPass4_frame_config bel_X3Y4_RES0 (.I0(W_RES0[23]), .I1(W_RES0[22]), .I2(W_RES0[21]), .I3(W_RES0[20]));
(* keep, BEL="X3Y4.OPB" *) InPass4_frame_config bel_X3Y4_OPB (.O0(W_OPB[23]), .O1(W_OPB[22]), .O2(W_OPB[21]), .O3(W_OPB[20]));
(* keep, BEL="X3Y4.OPA" *) InPass4_frame_config bel_X3Y4_OPA (.O0(W_OPA[23]), .O1(W_OPA[22]), .O2(W_OPA[21]), .O3(W_OPA[20]));
(* keep, BEL="X3Y3.RES2" *) OutPass4_frame_config bel_X3Y3_RES2 (.I0(W_RES2[27]), .I1(W_RES2[26]), .I2(W_RES2[25]), .I3(W_RES2[24]));
(* keep, BEL="X3Y3.RES1" *) OutPass4_frame_config bel_X3Y3_RES1 (.I0(W_RES1[27]), .I1(W_RES1[26]), .I2(W_RES1[25]), .I3(W_RES1[24]));
(* keep, BEL="X3Y3.RES0" *) OutPass4_frame_config bel_X3Y3_RES0 (.I0(W_RES0[27]), .I1(W_RES0[26]), .I2(W_RES0[25]), .I3(W_RES0[24]));
(* keep, BEL="X3Y3.OPB" *) InPass4_frame_config bel_X3Y3_OPB (.O0(W_OPB[27]), .O1(W_OPB[26]), .O2(W_OPB[25]), .O3(W_OPB[24]));
(* keep, BEL="X3Y3.OPA" *) InPass4_frame_config bel_X3Y3_OPA (.O0(W_OPA[27]), .O1(W_OPA[26]), .O2(W_OPA[25]), .O3(W_OPA[24]));
(* keep, BEL="X3Y2.RES2" *) OutPass4_frame_config bel_X3Y2_RES2 (.I0(W_RES2[31]), .I1(W_RES2[30]), .I2(W_RES2[29]), .I3(W_RES2[28]));
(* keep, BEL="X3Y2.RES1" *) OutPass4_frame_config bel_X3Y2_RES1 (.I0(W_RES1[31]), .I1(W_RES1[30]), .I2(W_RES1[29]), .I3(W_RES1[28]));
(* keep, BEL="X3Y2.RES0" *) OutPass4_frame_config bel_X3Y2_RES0 (.I0(W_RES0[31]), .I1(W_RES0[30]), .I2(W_RES0[29]), .I3(W_RES0[28]));
(* keep, BEL="X3Y2.OPB" *) InPass4_frame_config bel_X3Y2_OPB (.O0(W_OPB[31]), .O1(W_OPB[30]), .O2(W_OPB[29]), .O3(W_OPB[28]));
(* keep, BEL="X3Y2.OPA" *) InPass4_frame_config bel_X3Y2_OPA (.O0(W_OPA[31]), .O1(W_OPA[30]), .O2(W_OPA[29]), .O3(W_OPA[28]));
(* keep, BEL="X3Y1.RES2" *) OutPass4_frame_config bel_X3Y1_RES2 (.I0(W_RES2[35]), .I1(W_RES2[34]), .I2(W_RES2[33]), .I3(W_RES2[32]));
(* keep, BEL="X3Y1.RES1" *) OutPass4_frame_config bel_X3Y1_RES1 (.I0(W_RES1[35]), .I1(W_RES1[34]), .I2(W_RES1[33]), .I3(W_RES1[32]));
(* keep, BEL="X3Y1.RES0" *) OutPass4_frame_config bel_X3Y1_RES0 (.I0(W_RES0[35]), .I1(W_RES0[34]), .I2(W_RES0[33]), .I3(W_RES0[32]));
(* keep, BEL="X3Y1.OPB" *) InPass4_frame_config bel_X3Y1_OPB (.O0(W_OPB[35]), .O1(W_OPB[34]), .O2(W_OPB[33]), .O3(W_OPB[32]));
(* keep, BEL="X3Y1.OPA" *) InPass4_frame_config bel_X3Y1_OPA (.O0(W_OPA[35]), .O1(W_OPA[34]), .O2(W_OPA[33]), .O3(W_OPA[32]));
(* keep, BEL="X11Y9.RES2" *) OutPass4_frame_config bel_X11Y9_RES2 (.I0(E_RES2[3]), .I1(E_RES2[2]), .I2(E_RES2[1]), .I3(E_RES2[0]));
(* keep, BEL="X11Y9.RES1" *) OutPass4_frame_config bel_X11Y9_RES1 (.I0(E_RES1[3]), .I1(E_RES1[2]), .I2(E_RES1[1]), .I3(E_RES1[0]));
(* keep, BEL="X11Y9.RES0" *) OutPass4_frame_config bel_X11Y9_RES0 (.I0(E_RES0[3]), .I1(E_RES0[2]), .I2(E_RES0[1]), .I3(E_RES0[0]));
(* keep, BEL="X11Y9.OPB" *) InPass4_frame_config bel_X11Y9_OPB (.O0(E_OPB[3]), .O1(E_OPB[2]), .O2(E_OPB[1]), .O3(E_OPB[0]));
(* keep, BEL="X11Y9.OPA" *) InPass4_frame_config bel_X11Y9_OPA (.O0(E_OPA[3]), .O1(E_OPA[2]), .O2(E_OPA[1]), .O3(E_OPA[0]));
(* keep, BEL="X11Y8.RES2" *) OutPass4_frame_config bel_X11Y8_RES2 (.I0(E_RES2[7]), .I1(E_RES2[6]), .I2(E_RES2[5]), .I3(E_RES2[4]));
(* keep, BEL="X11Y8.RES1" *) OutPass4_frame_config bel_X11Y8_RES1 (.I0(E_RES1[7]), .I1(E_RES1[6]), .I2(E_RES1[5]), .I3(E_RES1[4]));
(* keep, BEL="X11Y8.RES0" *) OutPass4_frame_config bel_X11Y8_RES0 (.I0(E_RES0[7]), .I1(E_RES0[6]), .I2(E_RES0[5]), .I3(E_RES0[4]));
(* keep, BEL="X11Y8.OPB" *) InPass4_frame_config bel_X11Y8_OPB (.O0(E_OPB[7]), .O1(E_OPB[6]), .O2(E_OPB[5]), .O3(E_OPB[4]));
(* keep, BEL="X11Y8.OPA" *) InPass4_frame_config bel_X11Y8_OPA (.O0(E_OPA[7]), .O1(E_OPA[6]), .O2(E_OPA[5]), .O3(E_OPA[4]));
(* keep, BEL="X11Y7.RES2" *) OutPass4_frame_config bel_X11Y7_RES2 (.I0(E_RES2[11]), .I1(E_RES2[10]), .I2(E_RES2[9]), .I3(E_RES2[8]));
(* keep, BEL="X11Y7.RES1" *) OutPass4_frame_config bel_X11Y7_RES1 (.I0(E_RES1[11]), .I1(E_RES1[10]), .I2(E_RES1[9]), .I3(E_RES1[8]));
(* keep, BEL="X11Y7.RES0" *) OutPass4_frame_config bel_X11Y7_RES0 (.I0(E_RES0[11]), .I1(E_RES0[10]), .I2(E_RES0[9]), .I3(E_RES0[8]));
(* keep, BEL="X11Y7.OPB" *) InPass4_frame_config bel_X11Y7_OPB (.O0(E_OPB[11]), .O1(E_OPB[10]), .O2(E_OPB[9]), .O3(E_OPB[8]));
(* keep, BEL="X11Y7.OPA" *) InPass4_frame_config bel_X11Y7_OPA (.O0(E_OPA[11]), .O1(E_OPA[10]), .O2(E_OPA[9]), .O3(E_OPA[8]));
(* keep, BEL="X11Y6.RES2" *) OutPass4_frame_config bel_X11Y6_RES2 (.I0(E_RES2[15]), .I1(E_RES2[14]), .I2(E_RES2[13]), .I3(E_RES2[12]));
(* keep, BEL="X11Y6.RES1" *) OutPass4_frame_config bel_X11Y6_RES1 (.I0(E_RES1[15]), .I1(E_RES1[14]), .I2(E_RES1[13]), .I3(E_RES1[12]));
(* keep, BEL="X11Y6.RES0" *) OutPass4_frame_config bel_X11Y6_RES0 (.I0(E_RES0[15]), .I1(E_RES0[14]), .I2(E_RES0[13]), .I3(E_RES0[12]));
(* keep, BEL="X11Y6.OPB" *) InPass4_frame_config bel_X11Y6_OPB (.O0(E_OPB[15]), .O1(E_OPB[14]), .O2(E_OPB[13]), .O3(E_OPB[12]));
(* keep, BEL="X11Y6.OPA" *) InPass4_frame_config bel_X11Y6_OPA (.O0(E_OPA[15]), .O1(E_OPA[14]), .O2(E_OPA[13]), .O3(E_OPA[12]));
(* keep, BEL="X11Y5.RES2" *) OutPass4_frame_config bel_X11Y5_RES2 (.I0(E_RES2[19]), .I1(E_RES2[18]), .I2(E_RES2[17]), .I3(E_RES2[16]));
(* keep, BEL="X11Y5.RES1" *) OutPass4_frame_config bel_X11Y5_RES1 (.I0(E_RES1[19]), .I1(E_RES1[18]), .I2(E_RES1[17]), .I3(E_RES1[16]));
(* keep, BEL="X11Y5.RES0" *) OutPass4_frame_config bel_X11Y5_RES0 (.I0(E_RES0[19]), .I1(E_RES0[18]), .I2(E_RES0[17]), .I3(E_RES0[16]));
(* keep, BEL="X11Y5.OPB" *) InPass4_frame_config bel_X11Y5_OPB (.O0(E_OPB[19]), .O1(E_OPB[18]), .O2(E_OPB[17]), .O3(E_OPB[16]));
(* keep, BEL="X11Y5.OPA" *) InPass4_frame_config bel_X11Y5_OPA (.O0(E_OPA[19]), .O1(E_OPA[18]), .O2(E_OPA[17]), .O3(E_OPA[16]));
(* keep, BEL="X11Y4.RES2" *) OutPass4_frame_config bel_X11Y4_RES2 (.I0(E_RES2[23]), .I1(E_RES2[22]), .I2(E_RES2[21]), .I3(E_RES2[20]));
(* keep, BEL="X11Y4.RES1" *) OutPass4_frame_config bel_X11Y4_RES1 (.I0(E_RES1[23]), .I1(E_RES1[22]), .I2(E_RES1[21]), .I3(E_RES1[20]));
(* keep, BEL="X11Y4.RES0" *) OutPass4_frame_config bel_X11Y4_RES0 (.I0(E_RES0[23]), .I1(E_RES0[22]), .I2(E_RES0[21]), .I3(E_RES0[20]));
(* keep, BEL="X11Y4.OPB" *) InPass4_frame_config bel_X11Y4_OPB (.O0(E_OPB[23]), .O1(E_OPB[22]), .O2(E_OPB[21]), .O3(E_OPB[20]));
(* keep, BEL="X11Y4.OPA" *) InPass4_frame_config bel_X11Y4_OPA (.O0(E_OPA[23]), .O1(E_OPA[22]), .O2(E_OPA[21]), .O3(E_OPA[20]));
(* keep, BEL="X11Y3.RES2" *) OutPass4_frame_config bel_X11Y3_RES2 (.I0(E_RES2[27]), .I1(E_RES2[26]), .I2(E_RES2[25]), .I3(E_RES2[24]));
(* keep, BEL="X11Y3.RES1" *) OutPass4_frame_config bel_X11Y3_RES1 (.I0(E_RES1[27]), .I1(E_RES1[26]), .I2(E_RES1[25]), .I3(E_RES1[24]));
(* keep, BEL="X11Y3.RES0" *) OutPass4_frame_config bel_X11Y3_RES0 (.I0(E_RES0[27]), .I1(E_RES0[26]), .I2(E_RES0[25]), .I3(E_RES0[24]));
(* keep, BEL="X11Y3.OPB" *) InPass4_frame_config bel_X11Y3_OPB (.O0(E_OPB[27]), .O1(E_OPB[26]), .O2(E_OPB[25]), .O3(E_OPB[24]));
(* keep, BEL="X11Y3.OPA" *) InPass4_frame_config bel_X11Y3_OPA (.O0(E_OPA[27]), .O1(E_OPA[26]), .O2(E_OPA[25]), .O3(E_OPA[24]));
(* keep, BEL="X11Y2.RES2" *) OutPass4_frame_config bel_X11Y2_RES2 (.I0(E_RES2[31]), .I1(E_RES2[30]), .I2(E_RES2[29]), .I3(E_RES2[28]));
(* keep, BEL="X11Y2.RES1" *) OutPass4_frame_config bel_X11Y2_RES1 (.I0(E_RES1[31]), .I1(E_RES1[30]), .I2(E_RES1[29]), .I3(E_RES1[28]));
(* keep, BEL="X11Y2.RES0" *) OutPass4_frame_config bel_X11Y2_RES0 (.I0(E_RES0[31]), .I1(E_RES0[30]), .I2(E_RES0[29]), .I3(E_RES0[28]));
(* keep, BEL="X11Y2.OPB" *) InPass4_frame_config bel_X11Y2_OPB (.O0(E_OPB[31]), .O1(E_OPB[30]), .O2(E_OPB[29]), .O3(E_OPB[28]));
(* keep, BEL="X11Y2.OPA" *) InPass4_frame_config bel_X11Y2_OPA (.O0(E_OPA[31]), .O1(E_OPA[30]), .O2(E_OPA[29]), .O3(E_OPA[28]));
(* keep, BEL="X11Y1.RES2" *) OutPass4_frame_config bel_X11Y1_RES2 (.I0(E_RES2[35]), .I1(E_RES2[34]), .I2(E_RES2[33]), .I3(E_RES2[32]));
(* keep, BEL="X11Y1.RES1" *) OutPass4_frame_config bel_X11Y1_RES1 (.I0(E_RES1[35]), .I1(E_RES1[34]), .I2(E_RES1[33]), .I3(E_RES1[32]));
(* keep, BEL="X11Y1.RES0" *) OutPass4_frame_config bel_X11Y1_RES0 (.I0(E_RES0[35]), .I1(E_RES0[34]), .I2(E_RES0[33]), .I3(E_RES0[32]));
(* keep, BEL="X11Y1.OPB" *) InPass4_frame_config bel_X11Y1_OPB (.O0(E_OPB[35]), .O1(E_OPB[34]), .O2(E_OPB[33]), .O3(E_OPB[32]));
(* keep, BEL="X11Y1.OPA" *) InPass4_frame_config bel_X11Y1_OPA (.O0(E_OPA[35]), .O1(E_OPA[34]), .O2(E_OPA[33]), .O3(E_OPA[32]));
//(* keep, BEL="X14Y14.L" *) Config_access bel_X14Y14_L ();
(* keep, BEL="X14Y14.FAB2RAM_C" *) OutPass4_frame_config bel_X14Y14_FAB2RAM_C (.I0(OutPass4_frame_config_I0[54]), .I1(OutPass4_frame_config_I1[54]), .I2(OutPass4_frame_config_I2[54]), .I3(OutPass4_frame_config_I3[54]));
(* keep, BEL="X14Y14.FAB2RAM_A1" *) OutPass4_frame_config bel_X14Y14_FAB2RAM_A1 (.I0(OutPass4_frame_config_I0[55]), .I1(OutPass4_frame_config_I1[55]), .I2(OutPass4_frame_config_I2[55]), .I3(OutPass4_frame_config_I3[55]));
(* keep, BEL="X14Y14.FAB2RAM_A0" *) OutPass4_frame_config bel_X14Y14_FAB2RAM_A0 (.I0(OutPass4_frame_config_I0[56]), .I1(OutPass4_frame_config_I1[56]), .I2(OutPass4_frame_config_I2[56]), .I3(OutPass4_frame_config_I3[56]));
(* keep, BEL="X14Y14.FAB2RAM_D3" *) OutPass4_frame_config bel_X14Y14_FAB2RAM_D3 (.I0(OutPass4_frame_config_I0[57]), .I1(OutPass4_frame_config_I1[57]), .I2(OutPass4_frame_config_I2[57]), .I3(OutPass4_frame_config_I3[57]));
(* keep, BEL="X14Y14.FAB2RAM_D2" *) OutPass4_frame_config bel_X14Y14_FAB2RAM_D2 (.I0(OutPass4_frame_config_I0[58]), .I1(OutPass4_frame_config_I1[58]), .I2(OutPass4_frame_config_I2[58]), .I3(OutPass4_frame_config_I3[58]));
(* keep, BEL="X14Y14.FAB2RAM_D1" *) OutPass4_frame_config bel_X14Y14_FAB2RAM_D1 (.I0(OutPass4_frame_config_I0[59]), .I1(OutPass4_frame_config_I1[59]), .I2(OutPass4_frame_config_I2[59]), .I3(OutPass4_frame_config_I3[59]));
(* keep, BEL="X14Y14.FAB2RAM_D0" *) OutPass4_frame_config bel_X14Y14_FAB2RAM_D0 (.I0(OutPass4_frame_config_I0[60]), .I1(OutPass4_frame_config_I1[60]), .I2(OutPass4_frame_config_I2[60]), .I3(OutPass4_frame_config_I3[60]));
(* keep, BEL="X14Y14.RAM2FAB_D3" *) InPass4_frame_config bel_X14Y14_RAM2FAB_D3 (.O0(InPass4_frame_config_O0[36]), .O1(InPass4_frame_config_O1[36]), .O2(InPass4_frame_config_O2[36]), .O3(InPass4_frame_config_O3[36]));
(* keep, BEL="X14Y14.RAM2FAB_D2" *) InPass4_frame_config bel_X14Y14_RAM2FAB_D2 (.O0(InPass4_frame_config_O0[37]), .O1(InPass4_frame_config_O1[37]), .O2(InPass4_frame_config_O2[37]), .O3(InPass4_frame_config_O3[37]));
(* keep, BEL="X14Y14.RAM2FAB_D1" *) InPass4_frame_config bel_X14Y14_RAM2FAB_D1 (.O0(InPass4_frame_config_O0[38]), .O1(InPass4_frame_config_O1[38]), .O2(InPass4_frame_config_O2[38]), .O3(InPass4_frame_config_O3[38]));
(* keep, BEL="X14Y14.RAM2FAB_D0" *) InPass4_frame_config bel_X14Y14_RAM2FAB_D0 (.O0(InPass4_frame_config_O0[39]), .O1(InPass4_frame_config_O1[39]), .O2(InPass4_frame_config_O2[39]), .O3(InPass4_frame_config_O3[39]));
//(* keep, BEL="X14Y13.L" *) Config_access bel_X14Y13_L ();
(* keep, BEL="X14Y13.FAB2RAM_C" *) OutPass4_frame_config bel_X14Y13_FAB2RAM_C (.I0(OutPass4_frame_config_I0[61]), .I1(OutPass4_frame_config_I1[61]), .I2(OutPass4_frame_config_I2[61]), .I3(OutPass4_frame_config_I3[61]));
(* keep, BEL="X14Y13.FAB2RAM_A1" *) OutPass4_frame_config bel_X14Y13_FAB2RAM_A1 (.I0(OutPass4_frame_config_I0[62]), .I1(OutPass4_frame_config_I1[62]), .I2(OutPass4_frame_config_I2[62]), .I3(OutPass4_frame_config_I3[62]));
(* keep, BEL="X14Y13.FAB2RAM_A0" *) OutPass4_frame_config bel_X14Y13_FAB2RAM_A0 (.I0(OutPass4_frame_config_I0[63]), .I1(OutPass4_frame_config_I1[63]), .I2(OutPass4_frame_config_I2[63]), .I3(OutPass4_frame_config_I3[63]));
(* keep, BEL="X14Y13.FAB2RAM_D3" *) OutPass4_frame_config bel_X14Y13_FAB2RAM_D3 (.I0(OutPass4_frame_config_I0[64]), .I1(OutPass4_frame_config_I1[64]), .I2(OutPass4_frame_config_I2[64]), .I3(OutPass4_frame_config_I3[64]));
(* keep, BEL="X14Y13.FAB2RAM_D2" *) OutPass4_frame_config bel_X14Y13_FAB2RAM_D2 (.I0(OutPass4_frame_config_I0[65]), .I1(OutPass4_frame_config_I1[65]), .I2(OutPass4_frame_config_I2[65]), .I3(OutPass4_frame_config_I3[65]));
(* keep, BEL="X14Y13.FAB2RAM_D1" *) OutPass4_frame_config bel_X14Y13_FAB2RAM_D1 (.I0(OutPass4_frame_config_I0[66]), .I1(OutPass4_frame_config_I1[66]), .I2(OutPass4_frame_config_I2[66]), .I3(OutPass4_frame_config_I3[66]));
(* keep, BEL="X14Y13.FAB2RAM_D0" *) OutPass4_frame_config bel_X14Y13_FAB2RAM_D0 (.I0(OutPass4_frame_config_I0[67]), .I1(OutPass4_frame_config_I1[67]), .I2(OutPass4_frame_config_I2[67]), .I3(OutPass4_frame_config_I3[67]));
(* keep, BEL="X14Y13.RAM2FAB_D3" *) InPass4_frame_config bel_X14Y13_RAM2FAB_D3 (.O0(InPass4_frame_config_O0[40]), .O1(InPass4_frame_config_O1[40]), .O2(InPass4_frame_config_O2[40]), .O3(InPass4_frame_config_O3[40]));
(* keep, BEL="X14Y13.RAM2FAB_D2" *) InPass4_frame_config bel_X14Y13_RAM2FAB_D2 (.O0(InPass4_frame_config_O0[41]), .O1(InPass4_frame_config_O1[41]), .O2(InPass4_frame_config_O2[41]), .O3(InPass4_frame_config_O3[41]));
(* keep, BEL="X14Y13.RAM2FAB_D1" *) InPass4_frame_config bel_X14Y13_RAM2FAB_D1 (.O0(InPass4_frame_config_O0[42]), .O1(InPass4_frame_config_O1[42]), .O2(InPass4_frame_config_O2[42]), .O3(InPass4_frame_config_O3[42]));
(* keep, BEL="X14Y13.RAM2FAB_D0" *) InPass4_frame_config bel_X14Y13_RAM2FAB_D0 (.O0(InPass4_frame_config_O0[43]), .O1(InPass4_frame_config_O1[43]), .O2(InPass4_frame_config_O2[43]), .O3(InPass4_frame_config_O3[43]));
//(* keep, BEL="X14Y12.L" *) Config_access bel_X14Y12_L ();
(* keep, BEL="X14Y12.FAB2RAM_C" *) OutPass4_frame_config bel_X14Y12_FAB2RAM_C (.I0(OutPass4_frame_config_I0[68]), .I1(OutPass4_frame_config_I1[68]), .I2(OutPass4_frame_config_I2[68]), .I3(OutPass4_frame_config_I3[68]));
(* keep, BEL="X14Y12.FAB2RAM_A1" *) OutPass4_frame_config bel_X14Y12_FAB2RAM_A1 (.I0(OutPass4_frame_config_I0[69]), .I1(OutPass4_frame_config_I1[69]), .I2(OutPass4_frame_config_I2[69]), .I3(OutPass4_frame_config_I3[69]));
(* keep, BEL="X14Y12.FAB2RAM_A0" *) OutPass4_frame_config bel_X14Y12_FAB2RAM_A0 (.I0(OutPass4_frame_config_I0[70]), .I1(OutPass4_frame_config_I1[70]), .I2(OutPass4_frame_config_I2[70]), .I3(OutPass4_frame_config_I3[70]));
(* keep, BEL="X14Y12.FAB2RAM_D3" *) OutPass4_frame_config bel_X14Y12_FAB2RAM_D3 (.I0(OutPass4_frame_config_I0[71]), .I1(OutPass4_frame_config_I1[71]), .I2(OutPass4_frame_config_I2[71]), .I3(OutPass4_frame_config_I3[71]));
(* keep, BEL="X14Y12.FAB2RAM_D2" *) OutPass4_frame_config bel_X14Y12_FAB2RAM_D2 (.I0(OutPass4_frame_config_I0[72]), .I1(OutPass4_frame_config_I1[72]), .I2(OutPass4_frame_config_I2[72]), .I3(OutPass4_frame_config_I3[72]));
(* keep, BEL="X14Y12.FAB2RAM_D1" *) OutPass4_frame_config bel_X14Y12_FAB2RAM_D1 (.I0(OutPass4_frame_config_I0[73]), .I1(OutPass4_frame_config_I1[73]), .I2(OutPass4_frame_config_I2[73]), .I3(OutPass4_frame_config_I3[73]));
(* keep, BEL="X14Y12.FAB2RAM_D0" *) OutPass4_frame_config bel_X14Y12_FAB2RAM_D0 (.I0(OutPass4_frame_config_I0[74]), .I1(OutPass4_frame_config_I1[74]), .I2(OutPass4_frame_config_I2[74]), .I3(OutPass4_frame_config_I3[74]));
(* keep, BEL="X14Y12.RAM2FAB_D3" *) InPass4_frame_config bel_X14Y12_RAM2FAB_D3 (.O0(InPass4_frame_config_O0[44]), .O1(InPass4_frame_config_O1[44]), .O2(InPass4_frame_config_O2[44]), .O3(InPass4_frame_config_O3[44]));
(* keep, BEL="X14Y12.RAM2FAB_D2" *) InPass4_frame_config bel_X14Y12_RAM2FAB_D2 (.O0(InPass4_frame_config_O0[45]), .O1(InPass4_frame_config_O1[45]), .O2(InPass4_frame_config_O2[45]), .O3(InPass4_frame_config_O3[45]));
(* keep, BEL="X14Y12.RAM2FAB_D1" *) InPass4_frame_config bel_X14Y12_RAM2FAB_D1 (.O0(InPass4_frame_config_O0[46]), .O1(InPass4_frame_config_O1[46]), .O2(InPass4_frame_config_O2[46]), .O3(InPass4_frame_config_O3[46]));
(* keep, BEL="X14Y12.RAM2FAB_D0" *) InPass4_frame_config bel_X14Y12_RAM2FAB_D0 (.O0(InPass4_frame_config_O0[47]), .O1(InPass4_frame_config_O1[47]), .O2(InPass4_frame_config_O2[47]), .O3(InPass4_frame_config_O3[47]));
//(* keep, BEL="X14Y11.L" *) Config_access bel_X14Y11_L ();
(* keep, BEL="X14Y11.FAB2RAM_C" *) OutPass4_frame_config bel_X14Y11_FAB2RAM_C (.I0(OutPass4_frame_config_I0[75]), .I1(OutPass4_frame_config_I1[75]), .I2(OutPass4_frame_config_I2[75]), .I3(OutPass4_frame_config_I3[75]));
(* keep, BEL="X14Y11.FAB2RAM_A1" *) OutPass4_frame_config bel_X14Y11_FAB2RAM_A1 (.I0(OutPass4_frame_config_I0[76]), .I1(OutPass4_frame_config_I1[76]), .I2(OutPass4_frame_config_I2[76]), .I3(OutPass4_frame_config_I3[76]));
(* keep, BEL="X14Y11.FAB2RAM_A0" *) OutPass4_frame_config bel_X14Y11_FAB2RAM_A0 (.I0(OutPass4_frame_config_I0[77]), .I1(OutPass4_frame_config_I1[77]), .I2(OutPass4_frame_config_I2[77]), .I3(OutPass4_frame_config_I3[77]));
(* keep, BEL="X14Y11.FAB2RAM_D3" *) OutPass4_frame_config bel_X14Y11_FAB2RAM_D3 (.I0(OutPass4_frame_config_I0[78]), .I1(OutPass4_frame_config_I1[78]), .I2(OutPass4_frame_config_I2[78]), .I3(OutPass4_frame_config_I3[78]));
(* keep, BEL="X14Y11.FAB2RAM_D2" *) OutPass4_frame_config bel_X14Y11_FAB2RAM_D2 (.I0(OutPass4_frame_config_I0[79]), .I1(OutPass4_frame_config_I1[79]), .I2(OutPass4_frame_config_I2[79]), .I3(OutPass4_frame_config_I3[79]));
(* keep, BEL="X14Y11.FAB2RAM_D1" *) OutPass4_frame_config bel_X14Y11_FAB2RAM_D1 (.I0(OutPass4_frame_config_I0[80]), .I1(OutPass4_frame_config_I1[80]), .I2(OutPass4_frame_config_I2[80]), .I3(OutPass4_frame_config_I3[80]));
(* keep, BEL="X14Y11.FAB2RAM_D0" *) OutPass4_frame_config bel_X14Y11_FAB2RAM_D0 (.I0(OutPass4_frame_config_I0[81]), .I1(OutPass4_frame_config_I1[81]), .I2(OutPass4_frame_config_I2[81]), .I3(OutPass4_frame_config_I3[81]));
(* keep, BEL="X14Y11.RAM2FAB_D3" *) InPass4_frame_config bel_X14Y11_RAM2FAB_D3 (.O0(InPass4_frame_config_O0[48]), .O1(InPass4_frame_config_O1[48]), .O2(InPass4_frame_config_O2[48]), .O3(InPass4_frame_config_O3[48]));
(* keep, BEL="X14Y11.RAM2FAB_D2" *) InPass4_frame_config bel_X14Y11_RAM2FAB_D2 (.O0(InPass4_frame_config_O0[49]), .O1(InPass4_frame_config_O1[49]), .O2(InPass4_frame_config_O2[49]), .O3(InPass4_frame_config_O3[49]));
(* keep, BEL="X14Y11.RAM2FAB_D1" *) InPass4_frame_config bel_X14Y11_RAM2FAB_D1 (.O0(InPass4_frame_config_O0[50]), .O1(InPass4_frame_config_O1[50]), .O2(InPass4_frame_config_O2[50]), .O3(InPass4_frame_config_O3[50]));
(* keep, BEL="X14Y11.RAM2FAB_D0" *) InPass4_frame_config bel_X14Y11_RAM2FAB_D0 (.O0(InPass4_frame_config_O0[51]), .O1(InPass4_frame_config_O1[51]), .O2(InPass4_frame_config_O2[51]), .O3(InPass4_frame_config_O3[51]));
//(* keep, BEL="X14Y10.L" *) Config_access bel_X14Y10_L ();
(* keep, BEL="X14Y10.FAB2RAM_C" *) OutPass4_frame_config bel_X14Y10_FAB2RAM_C (.I0(OutPass4_frame_config_I0[82]), .I1(OutPass4_frame_config_I1[82]), .I2(OutPass4_frame_config_I2[82]), .I3(OutPass4_frame_config_I3[82]));
(* keep, BEL="X14Y10.FAB2RAM_A1" *) OutPass4_frame_config bel_X14Y10_FAB2RAM_A1 (.I0(OutPass4_frame_config_I0[83]), .I1(OutPass4_frame_config_I1[83]), .I2(OutPass4_frame_config_I2[83]), .I3(OutPass4_frame_config_I3[83]));
(* keep, BEL="X14Y10.FAB2RAM_A0" *) OutPass4_frame_config bel_X14Y10_FAB2RAM_A0 (.I0(OutPass4_frame_config_I0[84]), .I1(OutPass4_frame_config_I1[84]), .I2(OutPass4_frame_config_I2[84]), .I3(OutPass4_frame_config_I3[84]));
(* keep, BEL="X14Y10.FAB2RAM_D3" *) OutPass4_frame_config bel_X14Y10_FAB2RAM_D3 (.I0(OutPass4_frame_config_I0[85]), .I1(OutPass4_frame_config_I1[85]), .I2(OutPass4_frame_config_I2[85]), .I3(OutPass4_frame_config_I3[85]));
(* keep, BEL="X14Y10.FAB2RAM_D2" *) OutPass4_frame_config bel_X14Y10_FAB2RAM_D2 (.I0(OutPass4_frame_config_I0[86]), .I1(OutPass4_frame_config_I1[86]), .I2(OutPass4_frame_config_I2[86]), .I3(OutPass4_frame_config_I3[86]));
(* keep, BEL="X14Y10.FAB2RAM_D1" *) OutPass4_frame_config bel_X14Y10_FAB2RAM_D1 (.I0(OutPass4_frame_config_I0[87]), .I1(OutPass4_frame_config_I1[87]), .I2(OutPass4_frame_config_I2[87]), .I3(OutPass4_frame_config_I3[87]));
(* keep, BEL="X14Y10.FAB2RAM_D0" *) OutPass4_frame_config bel_X14Y10_FAB2RAM_D0 (.I0(OutPass4_frame_config_I0[88]), .I1(OutPass4_frame_config_I1[88]), .I2(OutPass4_frame_config_I2[88]), .I3(OutPass4_frame_config_I3[88]));
(* keep, BEL="X14Y10.RAM2FAB_D3" *) InPass4_frame_config bel_X14Y10_RAM2FAB_D3 (.O0(InPass4_frame_config_O0[52]), .O1(InPass4_frame_config_O1[52]), .O2(InPass4_frame_config_O2[52]), .O3(InPass4_frame_config_O3[52]));
(* keep, BEL="X14Y10.RAM2FAB_D2" *) InPass4_frame_config bel_X14Y10_RAM2FAB_D2 (.O0(InPass4_frame_config_O0[53]), .O1(InPass4_frame_config_O1[53]), .O2(InPass4_frame_config_O2[53]), .O3(InPass4_frame_config_O3[53]));
(* keep, BEL="X14Y10.RAM2FAB_D1" *) InPass4_frame_config bel_X14Y10_RAM2FAB_D1 (.O0(InPass4_frame_config_O0[54]), .O1(InPass4_frame_config_O1[54]), .O2(InPass4_frame_config_O2[54]), .O3(InPass4_frame_config_O3[54]));
(* keep, BEL="X14Y10.RAM2FAB_D0" *) InPass4_frame_config bel_X14Y10_RAM2FAB_D0 (.O0(InPass4_frame_config_O0[55]), .O1(InPass4_frame_config_O1[55]), .O2(InPass4_frame_config_O2[55]), .O3(InPass4_frame_config_O3[55]));


// bel IO_1_bidirectional_frame_config_pass input wires:
wire [9:0]IO_1_bidirectional_frame_config_pass_I;
wire [9:0]IO_1_bidirectional_frame_config_pass_T;
// bel IO_1_bidirectional_frame_config_pass output wires:
wire [9:0]IO_1_bidirectional_frame_config_pass_O;
wire [9:0]IO_1_bidirectional_frame_config_pass_Q;
// bel OutPass4_frame_config input wires:
wire [88:0]OutPass4_frame_config_I0;
wire [88:0]OutPass4_frame_config_I1;
wire [88:0]OutPass4_frame_config_I2;
wire [88:0]OutPass4_frame_config_I3;
// bel InPass4_frame_config output wires:
wire [55:0]InPass4_frame_config_O0;
wire [55:0]InPass4_frame_config_O1;
wire [55:0]InPass4_frame_config_O2;
wire [55:0]InPass4_frame_config_O3;

wire [35:0] W_OPA;
wire [35:0] W_OPB;
wire [35:0] W_RES0;
wire [35:0] W_RES1;
wire [35:0] W_RES2;
wire [35:0] E_OPA;
wire [35:0] E_OPB;
wire [35:0] E_RES0;
wire [35:0] E_RES1;
wire [35:0] E_RES2;

// instantiate user_design
top user_design_i (
    .clk(clk),
    .W_OPA(W_OPA),
    .W_OPB(W_OPB),
    .W_RES0(W_RES0),
    .W_RES1(W_RES1),
    .W_RES2(W_RES2),
    .E_OPA(E_OPA),
    .E_OPB(E_OPB),
    .E_RES0(E_RES0),
    .E_RES1(E_RES1),
    .E_RES2(E_RES2),
    .io_in(IO_1_bidirectional_frame_config_pass_O),
    .io_out(IO_1_bidirectional_frame_config_pass_I),
    .io_oeb(IO_1_bidirectional_frame_config_pass_T)
);


endmodule //top_wrapper
